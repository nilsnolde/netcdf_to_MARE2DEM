netcdf STOS_01Tx002a_01Rx001a_rotated {
dimensions:
	nx = 1 ;
	ny = 1 ;
	nz = 1 ;
	nogrid = 1 ;
	nsamp = UNLIMITED ; // (6360 currently)
	jtrace = 1 ;
	strace = 6 ;
	j_noisetrace = 1 ;
	j_masktrace = 1 ;
	csamp = 318 ;
	ttrace = 2 ;
	dtrace = 4 ;
	d_noisetrace = 4 ;
	d_masktrace = 4 ;
variables:
	float grid(nx, ny, nz, nogrid) ;
		grid:grid_trace = 0 ;
		grid:grid_fieldtype = "none" ;
		grid:grid_dx = 0.f ;
		grid:grid_dy = 0.f ;
		grid:grid_dz = 0.f ;
		grid:grid_x0 = 0.f ;
		grid:grid_y0 = 0.f ;
		grid:grid_z0 = 0.f ;
		grid:grid_undefined = -1.f ;
	float jsrc(nsamp, jtrace) ;
		jsrc:jsrc_trace = 1 ;
		jsrc:jsrc_fieldtype = "Jx" ;
		jsrc:jsrc_units = "A" ;
		jsrc:jsrc_undefined = -1.f ;
	float srcpos(nsamp, strace) ;
		srcpos:srcpos_trace = 6 ;
		srcpos:srcpos_direction = "x y z wd hd _" ;
		srcpos:srcpos_units = "m m m m deg _" ;
		srcpos:srcpos_undefined = -1.f ;
	float jsrc_noise(nsamp, j_noisetrace) ;
		jsrc_noise:jsrc_trace = 1 ;
		jsrc_noise:jsrc_fieldtype = "Jx" ;
	float jsrc_mask(nsamp, j_masktrace) ;
		jsrc_mask:jsrc_trace = 1 ;
		jsrc_mask:jsrc_fieldtype = "Jx" ;
	float sigma_c(csamp) ;
		sigma_c:sigma_c_trace = 1 ;
		sigma_c:sigma_c_dt = 0.f ;
	double time(nsamp, ttrace) ;
		time:time_trace = 2 ;
		time:time_fieldtype = "start stop" ;
	float emf(nsamp, dtrace) ;
		emf:emf_trace = 4 ;
		emf:emf_fieldtype = "Ex Ey Hx Hy" ;
		emf:emf_calstat = "emgs-E00420208 emgs-E00421973 mfs8u0412 mfs8u0428" ;
		emf:emf_sign = 1, 1, 1, 1 ;
		emf:emf_gain = 1.f, 1.f, 1.f, 1.f ;
		emf:emf_scalefactor = 1.f, 1.f, 1.f, 1.f ;
		emf:emf_quality = 2, 2, 2, 2 ;
		emf:emf_dcvalue = 0.f, 0.f, 0.f, 0.f ;
		emf:emf_armlength = 7.98f, 7.98f, 0.f, 0.f ;
		emf:emf_transform_number = 1, 1, 1, 1 ;
		emf:emf_gain_type = "auto_gain auto_gain auto_gain auto_gain" ;
		emf:emf_undefined = -1.f ;
		emf:emf_units = "V/Am^2 V/Am^2 1/m^2 1/m^2" ;
	float emf_noise(nsamp, d_noisetrace) ;
		emf_noise:emf_trace = 4 ;
		emf_noise:emf_fieldtype = "Ex Ey Hx Hy" ;
	float emf_mask(nsamp, d_masktrace) ;
		emf_mask:emf_trace = 4 ;
		emf_mask:emf_fieldtype = "Ex Ey Hx Hy" ;

// global attributes:
		:version = "1.1.0" ;
		:prochist = "/home/oh/SBLwiz_v1.20.13969_emgs/bin/elsource2h5_R-1-8-0 innav=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/RawData/Navigation inawl=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/SurveyPlan/EMGS_8960ms_1357_80ms_squarewave.awl incrs=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/NavArchive/SBL_OnlineData/tx_P294 sourceNavRegular=on sourceCurrDownSampFactor=1 insource=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/.AntFiles/Source ofelmask=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/Source/?.h5src client=ShellTodd_NewZealand survey_area=Tasman_Sea vessel=Galatea survey_date=Jan_Feb_2011 source=01Tx002 freqs=0.111607142857,0.334821428571,0.558035714286,0.78125,1.00446428571,1.22767857143,1.45089285714,1.67410714286,1.89732142857,2.12053571429 verbose=5 logfile=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/SourceLogs/01Tx002.log ;/home/oh/SBLwiz_v1.20.0.13996_emgs_vessel/bin/elise_R-6-2-0 nred.fff_remove=on rawoutput=off channels=all rsamp=on temperature=4.00 ecal.armlen.z=2.00 ecal.armlen.y=7.98 ecal.armlen.x=7.98 gse.minGainLen=120 nred.flasherase.Jun08=eh ecal.impcomp.rmax=30.00 nred.despike.Dec06.std.e=8.00 gse.predLen=10 hcal.crosstalk_remove=on nred.despike.Dec06.std.h=8.00 ecal.impcomp=on ecal=on nred.despike.Dec06=eh elisefilterdir=/project/elmap/share/elisefilters/50Hz gse.flow=0.05 nred.flasherase.Jun08.length=500 hcal=on ifel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/RawData/Receiver/01Rx001a/STOS_01Rx001a_040211_061022.bin ofel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/Receivers/STOS_01Rx001a.h5 ofel2=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/DownsampledReceivers/STOS_01Rx001a.h5qc ofel2.downsample=50 logfile=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/ReceiverLogs/STOS_01Rx001a.txt verbose=5 ;/home/oh/SBLwiz_v1.20.0.13996_emgs_vessel/bin/elsetrecnav_R-1-6-0 vessel=Galatea survey_area=Tasman_Sea client=ShellTodd_NewZealand survey_date=Jan_Feb_2011 author=Oystein_Hallanger-Martin_Hansen innav=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/RawData/Navigation incrs=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/RawData/../NavArchive/SBL_OnlineData iofel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/Receivers/STOS_01Rx001a.h5 ;/home/mhansen/SBLwiz_v1.20.0.13996_emgs/bin/elsetrecnav_R-1-6 vessel=Galatea survey_area=Tasman_Sea client=ShellTodd_NewZealand survey_date=Jan_Feb_2011 author=Oystein_Hallanger-Martin_Hansen innav=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/RawData/Navigation incrs=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/RawData/../NavArchive/SBL_OnlineData iofel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/Receivers/STOS_01Rx001a.h5 ;/home/mhansen/SBLwiz_v1.20.0.13996_emgs/bin/eldemod_R-9-6-1 exclude_dc_noisegate=true zeropadding=off avgsp=on npmax=18 avgsr=on sn_separation_f=0.022321429 npmin=18 wintype=hanning mode=LINEOFFSET signal_gate_f=0.0 stoptime=2011-01-17-21:35:13 snr=on windowposmethod=ZEROOFFSET noise_gate_f=0.0390625 exclude=46750,46760 npzof=18 dr=80 rmin=499 r0=-15000 rlow=500 rf=15000 compsensimp=on starttime=2011-01-17-08:35:43 rhigh=10000 towlinemask=01Tx002a sourcepath=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/Source inrec=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_CSEM/Receivers/STOS_01Rx001a.h5 ofel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_01Tx002a_re/Demod/STOS_01Tx002a_01Rx001a_demod.nc ;/home/mhansen/SBLwiz_v1.20.0.13996_emgs/bin/elscale_R-1-3 mode=none2magphase ifel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_01Tx002a_re/Demod/STOS_01Tx002a_01Rx001a_demod.nc ofel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_01Tx002a_re/Scaled/STOS_01Tx002a_01Rx001a_scaled.nc ;/home/mhansen/SBLwiz_v1.20.0.13996_emgs/bin/eladd_R-4-0 saturated_window=2000 ey1=near ey2=far ex2=far ex1=all ifel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_01Tx002a_re/Scaled/STOS_01Tx002a_01Rx001a_scaled.nc ofel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_01Tx002a_re/Summed/STOS_01Tx002a_01Rx001a_summed.nc ;/home/mhansen/SBLwiz_v1.20.0.13996_emgs/bin/elrotate_R-3-0 angle_uncertainty=3.0 angle=261.269582 recheading=305.530000 ifel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_01Tx002a_re/Summed/STOS_01Tx002a_01Rx001a_summed.nc ofel=/mnt/ibrix3/surveys/Shell_Todd_New_Zealand/2011_Galatea/STOS/04_GSO_Reprocessing_May2011/Job_01Tx002a_re/Rotated/STOS_01Tx002a_01Rx001a_rotated.nc ;" ;
		:loghist = "elsource2h5 - $Name: R-1-8 $ $Date: 2011-20-04 15:44:56 $;Elise - $Name: R-6-2 $ $Date: 2011-04-17 15:44:56 $;elsetrecnav - $Name: R-1-6 $ $Date: 2011-04-10 15:44:56 $;elsetrecnav - $Name: R-1-6 $ $Date: 2011-04-10 15:44:56 $;eldemod - $Version: R-9-6-1 $ $Date: 2008-01-09 19:08:04 $;elscale - $Version: R-1-3 $ $Date: 2008-01-07 08:58:13 $;eladd - $Version: R-4-0 $ $Date: 2008-01-07 08:58:13 $;elrotate - Name: R-3-0;" ;
		:logid = "unknown" ;
		:surveyid = "STOS" ;
		:jobid = "unknown" ;
		:recid = "01Rx001a" ;
		:lineid = "01Tx002a" ;
		:domain = "frequency" ;
		:coilid = "unknown" ;
		:x_r = 1633491.f ;
		:y_r = 5619388.f ;
		:z_r = 109.4f ;
		:psi = 0.f ;
		:phi = 44.26042f ;
		:theta = 0.f ;
		:psi_uncertainty = 0.f ;
		:phi_uncertainty = 3.f ;
		:theta_uncertainty = 0.f ;
		:receiver_heading = -1000.f ;
		:sigma_f = 0.f ;
		:dataset_date = "Jan Feb 2011" ;
		:dataset_author = "Oystein Hallanger-Martin Hansen" ;
		:dlength = 270.52f ;
		:geodetic_datum = "unknown" ;
		:projection_type = "transverse_mercator_north_oriented" ;
		:projection_zone = "unknown" ;
		:long_of_central_meridian = "173deg 00min 00.000sec E" ;
		:grid_origin = "000deg 00min 00.000sec N,   173deg 00min 00.000sec E" ;
		:grid_coord_at_origin = "1600000.00E,  10000000.00N" ;
		:scale_factor = "unknown" ;
		:scale_factor_long_lat = "0.99960000000000004" ;
		:planned_vessel_speed = "2.00 kts" ;
		:format_type = "complex_demod" ;
		:t0_emgs = "17-01-2011 08:35:43" ;
		:t0_unix = 1295253343. ;
		:nf = 10 ;
		:freqs = 0.1116071f, 0.3348214f, 0.5580357f, 0.78125f, 1.004464f, 1.227679f, 1.450893f, 1.674107f, 1.897321f, 2.120536f ;
		:dx1 = 0.f ;
		:dx2 = 0.f ;
		:dk1 = 0.f ;
		:dk2 = 0.f ;
		:dt = 0.02f ;
		:clock_drift_ppb = 58.06309f ;
		:approx_source_heading = 44.26042f ;
data:

 grid =
  _ ;

 jsrc =
  851.5497,
  1334.176,
  851.7628,
  1333.763,
  850.7783,
  1334.407,
  851.3549,
  1334.604,
  851.6039,
  1334.059,
  852.0295,
  1334.351,
  851.5128,
  1334.632,
  851.7574,
  1334.235,
  851.6926,
  1334.123,
  852.2081,
  1333.977,
  851.5474,
  1333.309,
  852.3996,
  1333.003,
  851.8854,
  1334.323,
  852.0712,
  1334.182,
  852.8131,
  1333.978,
  851.8556,
  1334.473,
  851.277,
  1334.323,
  851.7197,
  1333.239,
  851.713,
  1333.394,
  851.1327,
  1332.731,
  850.1468,
  1331.851,
  850.8623,
  1332.388,
  850.6614,
  1334.117,
  851.5204,
  1334.42,
  851.8162,
  1333.42,
  851.4053,
  1333.456,
  851.6202,
  1333.489,
  851.5677,
  1333.806,
  852.425,
  1332.986,
  851.3555,
  1333.457,
  851.9053,
  1333.692,
  852.9982,
  1334.12,
  852.447,
  1334.268,
  851.7476,
  1334.673,
  852.1924,
  1334.084,
  852.2639,
  1334.124,
  851.1191,
  1334.585,
  851.5846,
  1334.264,
  851.9114,
  1334.509,
  851.6002,
  1334.868,
  851.5359,
  1334.665,
  851.6472,
  1334.824,
  851.8442,
  1334.157,
  852.3253,
  1333.805,
  852.6849,
  1333.324,
  852.1635,
  1333.055,
  852.0715,
  1334.553,
  852.2643,
  1334.283,
  852.5503,
  1333.073,
  852.6456,
  1333,
  851.3979,
  1333.529,
  852.0196,
  1333.638,
  852.5549,
  1333.577,
  852.5194,
  1333.656,
  850.8351,
  1333.691,
  851.7248,
  1334.038,
  852.2759,
  1334.087,
  851.6208,
  1334.444,
  851.4178,
  1333.702,
  851.5169,
  1333.733,
  851.6017,
  1333.79,
  851.8281,
  1333.813,
  852.1267,
  1333.833,
  851.4827,
  1333.701,
  851.7807,
  1333.788,
  852.2953,
  1333.746,
  852.8468,
  1333.933,
  852.7632,
  1333.888,
  851.9421,
  1333.54,
  852.2387,
  1333.676,
  852.6745,
  1333.024,
  852.6483,
  1333.875,
  851.6016,
  1334.5,
  852.1445,
  1333.759,
  852.6953,
  1333.43,
  851.542,
  1333.604,
  851.3511,
  1333.831,
  851.9049,
  1333.792,
  852.4985,
  1333.804,
  851.8414,
  1334.428,
  851.7168,
  1334.567,
  851.6736,
  1333.705,
  851.9373,
  1333.523,
  851.9376,
  1333.678,
  851.4035,
  1334.328,
  851.5768,
  1333.936,
  851.6242,
  1334.079,
  852.0628,
  1333.395,
  852.476,
  1333.468,
  851.9061,
  1334.202,
  852.3094,
  1334.549,
  852.3283,
  1333.931,
  852.8773,
  1333.266,
  852.5342,
  1334.155,
  852.0713,
  1334.067,
  852.5269,
  1333.906,
  853.0667,
  1333.413,
  852.0969,
  1333.182,
  851.5302,
  1333.597,
  851.9824,
  1333.517,
  852.4921,
  1333.238,
  852.1439,
  1333.654,
  851.2886,
  1334.336,
  852.0663,
  1334.466,
  852.29,
  1333.829,
  851.2794,
  1333.954,
  850.2858,
  1333.238,
  851.2414,
  1333.376,
  851.9474,
  1333.009,
  851.884,
  1332.969,
  851.0743,
  1333.865,
  850.7581,
  1332.666,
  851.3239,
  1333.595,
  851.699,
  1333.525,
  851.5251,
  1333.28,
  851.2835,
  1333.909,
  851.8604,
  1333.873,
  852.0001,
  1333.268,
  852.6165,
  1333.097,
  851.8604,
  1333.151,
  851.5886,
  1333.363,
  851.7534,
  1333.471,
  852.5248,
  1332.733,
  852.6897,
  1332.675,
  851.9888,
  1333.38,
  852.0652,
  1333.658,
  852.4432,
  1333.392,
  852.5782,
  1333.402,
  851.8558,
  1334.152,
  851.8359,
  1334.196,
  852.3427,
  1333.713,
  852.6059,
  1332.679,
  851.4338,
  1333.287,
  851.5585,
  1334.157,
  851.7852,
  1333.009,
  852.7489,
  1333.331,
  852.0795,
  1334.066,
  851.1039,
  1333.816,
  851.7707,
  1333.904,
  852.5911,
  1333.7,
  851.7953,
  1334.108,
  851.4171,
  1334.386,
  851.6165,
  1333.918,
  851.9572,
  1333.581,
  850.9366,
  1333.806,
  850.8959,
  1333.819,
  851.3425,
  1333.727,
  851.5311,
  1333.24,
  852.0074,
  1332.969,
  851.8005,
  1333.347,
  851.2159,
  1333.208,
  851.9484,
  1333.802,
  852.1081,
  1333.939,
  852.5615,
  1334.003,
  851.9926,
  1333.613,
  851.4056,
  1333.601,
  852.1622,
  1333.292,
  852.6049,
  1333.268,
  852.8779,
  1333.183,
  852.0281,
  1333.755,
  852.0283,
  1333.986,
  852.3099,
  1333.224,
  852.9721,
  1333.387,
  852.0107,
  1333.946,
  851.6138,
  1333.612,
  851.7869,
  1332.771,
  852.4282,
  1332.972,
  851.5849,
  1333.74,
  851.3332,
  1334.225,
  851.9309,
  1333.168,
  852.5082,
  1333.198,
  851.2383,
  1333.366,
  851.4672,
  1334.076,
  851.7676,
  1333.335,
  852.0742,
  1333.672,
  851.407,
  1334.648,
  851.2115,
  1334.278,
  851.6981,
  1334.298,
  852.153,
  1333.626,
  852.2222,
  1333.829,
  850.9917,
  1334.007,
  851.1597,
  1333.674,
  851.6719,
  1333.273,
  852.0623,
  1333.617,
  851.605,
  1334.177,
  851.1852,
  1334.144,
  851.7872,
  1333.526,
  852.2977,
  1333.406,
  852.2408,
  1333.261,
  851.6871,
  1334.018,
  851.3952,
  1334.114,
  852.1069,
  1333.951,
  852.6785,
  1333.392,
  852.5118,
  1334.194,
  851.6865,
  1334.318,
  851.6381,
  1333.26,
  852.2893,
  1333.281,
  852.2809,
  1333.151,
  852.6695,
  1333.619,
  851.9109,
  1333.672,
  852.0106,
  1333.158,
  852.6472,
  1332.949,
  853.0255,
  1333.491,
  851.877,
  1334.154,
  852.4498,
  1333.791,
  852.6179,
  1333.253,
  852.8058,
  1333.65,
  851.7786,
  1334.064,
  851.6938,
  1333.955,
  851.9334,
  1333.511,
  852.4033,
  1333.061,
  850.5536,
  1332.839,
  850.6955,
  1332.58,
  851.3956,
  1332.426,
  852.4336,
  1333.734,
  851.2337,
  1334.54,
  851.9149,
  1334.505,
  852.1384,
  1334.092,
  851.2134,
  1331.698,
  850.5117,
  1332.724,
  851.0878,
  1333.646,
  851.0742,
  1332.476,
  851.435,
  1331.762,
  851.9213,
  1333.158,
  851.3976,
  1334.448,
  851.6369,
  1333.902,
  851.4257,
  1332.621,
  851.048,
  1331.617,
  850.4487,
  1331.618,
  850.5449,
  1332.828,
  851.4195,
  1333.225,
  852.0104,
  1333.377,
  852.0234,
  1333.806,
  851.2239,
  1333.723,
  851.3857,
  1332.535,
  852.0268,
  1332.709,
  851.6884,
  1332.044,
  851.4749,
  1333.288,
  851.5435,
  1333.118,
  851.942,
  1333.513,
  852.2932,
  1333.15,
  852.4493,
  1333.866,
  852.1677,
  1334.006,
  851.9882,
  1333.736,
  852.1757,
  1333.391,
  851.9545,
  1332.254,
  851.0631,
  1332.935,
  851.0143,
  1333.151,
  851.7201,
  1333.435,
  852.5787,
  1333.554,
  852.9131,
  1333.638,
  851.4594,
  1333.34,
  851.7991,
  1333.229,
  851.954,
  1332.742,
  852.1061,
  1332.402,
  851.8633,
  1334.635,
  851.4067,
  1333.633,
  851.9152,
  1333.162,
  852.4062,
  1333.455,
  850.9556,
  1333.546,
  851.1171,
  1333.792,
  852.205,
  1334.102,
  852.8145,
  1334.384,
  852.0862,
  1334.488,
  850.9319,
  1333.814,
  850.9888,
  1332.499,
  852.0356,
  1332.992,
  851.7101,
  1334.147,
  851.485,
  1334.173,
  851.8638,
  1333.884,
  851.778,
  1333.458,
  851.9166,
  1333.93,
  851.4718,
  1334.465,
  851.6027,
  1334.693,
  851.4721,
  1333.774,
  852.4203,
  1333.409,
  851.547,
  1334.342,
  851.6064,
  1334.6,
  852.2032,
  1333.349,
  852.0383,
  1332.961,
  852.6186,
  1333.843,
  851.8724,
  1334.049,
  851.701,
  1334.122,
  852.0712,
  1333.534,
  852.5389,
  1333.596,
  852.1265,
  1333.442,
  851.7627,
  1333.527,
  851.6763,
  1333.593,
  852.0119,
  1333.438,
  852.2369,
  1332.86,
  852.5193,
  1334.273,
  851.9229,
  1333.975,
  852.108,
  1333.771,
  852.3723,
  1333.63,
  852.3516,
  1333.84,
  851.9553,
  1334.098,
  851.8051,
  1333.563,
  852.6718,
  1333.983,
  852.5692,
  1333.211,
  851.8157,
  1334.455,
  851.5619,
  1334.044,
  852.3262,
  1333.919,
  852.7068,
  1333.23,
  852.126,
  1334.134,
  851.8212,
  1334.683,
  852.5853,
  1334.516,
  852.1899,
  1333.129,
  851.3905,
  1333.859,
  851.362,
  1334.362,
  851.9443,
  1334.132,
  852.599,
  1334.072,
  851.8901,
  1334.418,
  851.3845,
  1334.638,
  851.9304,
  1334.697,
  851.9725,
  1333.719,
  851.6259,
  1333.222,
  851.0075,
  1333.905,
  851.7493,
  1334.625,
  519.7802,
  -64.28521,
  519.6546,
  -64.66864,
  519.6701,
  -63.41517,
  519.8539,
  -63.842,
  519.6025,
  -64.48195,
  519.8022,
  -64.73811,
  519.8862,
  -64.03316,
  519.8618,
  -64.53721,
  519.7672,
  -64.30668,
  519.8412,
  -64.98522,
  519.2916,
  -64.62182,
  519.3942,
  -65.30912,
  519.8595,
  -64.54221,
  519.8901,
  -64.71459,
  519.8154,
  -65.41842,
  519.8392,
  -64.34736,
  519.675,
  -64.07482,
  519.5275,
  -64.80467,
  519.3763,
  -64.80488,
  519.2479,
  -64.59169,
  518.5397,
  -64.40399,
  518.9365,
  -64.56287,
  519.4427,
  -63.76083,
  519.6937,
  -64.30432,
  519.3564,
  -64.86456,
  519.4211,
  -64.86903,
  519.5379,
  -64.78953,
  519.5488,
  -64.54357,
  519.434,
  -65.70343,
  519.5198,
  -64.1963,
  519.634,
  -64.89812,
  519.8252,
  -65.51267,
  519.8546,
  -64.91907,
  519.8517,
  -64.17598,
  519.907,
  -64.91131,
  519.6384,
  -64.86545,
  519.6287,
  -63.7171,
  519.7628,
  -64.13966,
  519.8553,
  -64.38509,
  519.8579,
  -63.88451,
  519.8165,
  -63.92456,
  520.0143,
  -64.00154,
  519.7037,
  -64.53625,
  519.6889,
  -64.9436,
  519.6561,
  -65.43903,
  519.4431,
  -65.15311,
  519.7784,
  -64.55721,
  519.8908,
  -64.79597,
  519.5911,
  -65.71061,
  519.4147,
  -65.53185,
  519.4458,
  -64.02268,
  519.5652,
  -64.86841,
  519.6648,
  -65.42633,
  519.5977,
  -65.20053,
  519.5623,
  -63.65678,
  519.8153,
  -64.30057,
  519.8165,
  -64.87191,
  519.723,
  -64.06203,
  519.6648,
  -64.4756,
  519.5314,
  -64.41013,
  519.6109,
  -64.47796,
  519.7434,
  -64.61076,
  519.7136,
  -64.99113,
  519.6154,
  -64.2502,
  519.6818,
  -64.62143,
  519.8068,
  -64.91441,
  519.8793,
  -65.30537,
  519.8202,
  -65.13473,
  519.5635,
  -64.52541,
  519.5995,
  -65.04187,
  519.4946,
  -65.73891,
  519.6456,
  -65.27362,
  519.7908,
  -64.13757,
  519.5517,
  -64.91679,
  519.7275,
  -65.46037,
  519.5765,
  -64.34696,
  519.535,
  -64.03576,
  519.8119,
  -64.70412,
  519.6951,
  -65.16233,
  519.739,
  -64.52135,
  519.7821,
  -64.10966,
  519.6428,
  -64.54873,
  519.6032,
  -64.95603,
  519.6224,
  -64.95654,
  519.6882,
  -63.99006,
  519.5891,
  -64.34233,
  519.4331,
  -64.41148,
  519.3677,
  -65.18776,
  519.5643,
  -65.22095,
  519.7322,
  -64.44492,
  519.9083,
  -64.76956,
  519.8033,
  -64.99768,
  519.7544,
  -65.74144,
  519.7823,
  -65.10925,
  519.7333,
  -64.73656,
  519.7772,
  -65.14008,
  519.7048,
  -65.9931,
  519.4538,
  -65.12003,
  519.5204,
  -64.42334,
  519.7379,
  -64.70975,
  519.6737,
  -65.48908,
  519.6423,
  -64.99223,
  519.5602,
  -64.14556,
  519.5836,
  -64.88762,
  519.7009,
  -65.29745,
  519.5546,
  -64.31815,
  519.3743,
  -63.71979,
  519.4335,
  -64.61935,
  519.2815,
  -65.15148,
  519.2932,
  -64.81239,
  519.3652,
  -64.08134,
  519.0314,
  -64.37772,
  519.2619,
  -64.75968,
  519.4149,
  -64.99511,
  519.3351,
  -64.87889,
  519.5189,
  -64.1451,
  519.6989,
  -64.74201,
  519.6334,
  -65.23111,
  519.2404,
  -65.76547,
  519.4161,
  -64.97382,
  519.5562,
  -64.66821,
  519.3792,
  -64.61378,
  519.3951,
  -65.78966,
  519.4492,
  -65.98011,
  519.4615,
  -65.27163,
  519.6588,
  -65.08557,
  519.5052,
  -65.46244,
  519.5891,
  -65.69721,
  519.6517,
  -64.4816,
  519.8487,
  -64.6898,
  519.717,
  -65.25816,
  519.5002,
  -65.76576,
  519.2051,
  -64.50723,
  519.6624,
  -64.33996,
  519.3002,
  -64.79549,
  519.5312,
  -65.61179,
  519.6697,
  -64.73849,
  519.3495,
  -63.97675,
  519.4888,
  -64.71867,
  519.6259,
  -65.24891,
  519.6483,
  -64.38308,
  519.8994,
  -64.19482,
  519.7873,
  -64.34406,
  519.5423,
  -64.9282,
  519.4064,
  -63.93113,
  519.3761,
  -63.90613,
  519.4441,
  -64.14398,
  519.5666,
  -64.87122,
  519.4445,
  -65.15163,
  519.6024,
  -64.61747,
  519.2726,
  -64.36635,
  519.5041,
  -64.92031,
  519.5461,
  -65.31551,
  519.8532,
  -65.47117,
  519.5615,
  -64.65985,
  519.3996,
  -64.47256,
  519.4205,
  -64.98801,
  519.386,
  -65.72988,
  519.4802,
  -66.21149,
  519.6744,
  -64.94713,
  519.6096,
  -64.84073,
  519.4857,
  -65.4603,
  519.4763,
  -65.991,
  519.4877,
  -64.71246,
  519.4479,
  -64.56097,
  519.207,
  -65.15979,
  519.4111,
  -65.72861,
  519.4402,
  -64.48747,
  519.663,
  -64.41446,
  519.5642,
  -65.148,
  519.4908,
  -65.61143,
  519.1857,
  -64.71532,
  519.521,
  -64.30328,
  519.5034,
  -64.69628,
  519.6464,
  -65.21543,
  519.91,
  -63.85099,
  519.6807,
  -63.81718,
  519.7567,
  -64.49311,
  519.5383,
  -65.00141,
  519.5974,
  -64.90575,
  519.378,
  -63.86211,
  519.3093,
  -63.94358,
  519.2316,
  -64.95712,
  519.6579,
  -65.31467,
  519.7494,
  -64.57188,
  519.6158,
  -64.15247,
  519.4277,
  -64.83072,
  519.3632,
  -65.40605,
  519.2557,
  -65.14503,
  519.6674,
  -64.59401,
  519.6108,
  -64.49847,
  519.683,
  -65.08818,
  519.7249,
  -65.38684,
  519.6995,
  -65.18202,
  519.8093,
  -64.29969,
  519.6298,
  -64.72351,
  519.6848,
  -65.15885,
  519.4795,
  -65.1748,
  519.6439,
  -65.33092,
  519.4922,
  -64.7554,
  519.3016,
  -65.36372,
  519.4746,
  -65.64501,
  519.7414,
  -65.74952,
  519.6988,
  -64.49063,
  519.7921,
  -65.09763,
  519.5648,
  -65.42919,
  519.5931,
  -65.56893,
  519.6761,
  -64.3959,
  519.6067,
  -64.58701,
  519.4716,
  -65.10822,
  519.1008,
  -65.58367,
  518.9952,
  -64.04258,
  519.1182,
  -64.5162,
  519.127,
  -65.03859,
  519.5718,
  -65.30177,
  519.6617,
  -63.89734,
  519.633,
  -64.23932,
  519.5454,
  -64.84467,
  518.8149,
  -65.35345,
  519.0786,
  -63.99197,
  519.4317,
  -64.11294,
  519.1652,
  -64.47636,
  519.0493,
  -65.16273,
  519.4692,
  -65.31672,
  519.579,
  -64.12459,
  519.5222,
  -64.52475,
  518.9025,
  -64.87633,
  519.0333,
  -65.13192,
  518.6634,
  -64.87079,
  518.9929,
  -64.06666,
  519.0051,
  -64.72387,
  519.2665,
  -64.99319,
  519.5461,
  -64.87727,
  519.52,
  -64.28239,
  519.1118,
  -64.96161,
  519.0757,
  -65.18427,
  519.011,
  -65.40358,
  519.407,
  -64.8838,
  519.2115,
  -64.74119,
  519.497,
  -65.01114,
  519.5109,
  -65.37376,
  519.8886,
  -65.07843,
  519.8279,
  -64.84489,
  519.5349,
  -64.77406,
  519.3699,
  -65.33438,
  518.9561,
  -65.80765,
  518.9268,
  -64.687,
  519.168,
  -64.3685,
  519.4934,
  -64.95905,
  519.639,
  -65.56664,
  519.5311,
  -65.76082,
  519.1941,
  -64.63395,
  519.3852,
  -64.66651,
  519.1432,
  -65.26411,
  518.8606,
  -65.69324,
  519.7087,
  -64.44773,
  519.5456,
  -64.4073,
  519.4763,
  -65.04738,
  519.6891,
  -65.4501,
  519.2885,
  -63.92937,
  519.4232,
  -64.08545,
  519.6456,
  -64.83118,
  519.7874,
  -65.26269,
  519.6841,
  -64.6958,
  519.3282,
  -63.99442,
  518.864,
  -64.48833,
  519.4149,
  -65.18848,
  519.623,
  -64.66851,
  519.769,
  -64.26911,
  519.7789,
  -64.78822,
  519.4631,
  -64.87582,
  519.556,
  -64.79758,
  519.4897,
  -64.09717,
  519.778,
  -63.99515,
  519.48,
  -64.45,
  519.4949,
  -65.3895,
  519.6622,
  -64.18909,
  519.9698,
  -64.13309,
  519.5684,
  -65.05582,
  519.1638,
  -65.16589,
  519.7028,
  -65.28419,
  519.597,
  -64.6824,
  519.8127,
  -64.30213,
  519.5604,
  -64.8028,
  519.7018,
  -65.30223,
  519.4879,
  -65.40703,
  519.3834,
  -65.04025,
  519.4743,
  -64.65274,
  519.5764,
  -65.34512,
  519.3295,
  -65.91901,
  519.931,
  -65.35584,
  519.7925,
  -64.8234,
  519.6993,
  -64.90598,
  519.7782,
  -65.36382,
  519.7933,
  -65.18515,
  519.8298,
  -64.79614,
  519.5497,
  -64.65611,
  519.7551,
  -65.35136,
  519.5038,
  -65.7621,
  519.8785,
  -64.56815,
  519.6054,
  -64.59915,
  519.7165,
  -64.9603,
  519.6195,
  -65.65733,
  519.7383,
  -64.65781,
  519.8711,
  -64.176,
  519.8923,
  -64.81945,
  519.5141,
  -65.32977,
  519.65,
  -64.28492,
  519.8008,
  -63.96609,
  519.7262,
  -64.51041,
  519.8004,
  -65.1963,
  519.7828,
  -64.50761,
  519.7635,
  -63.89323,
  519.8181,
  -64.45503,
  519.5321,
  -64.99551,
  519.35,
  -64.98746,
  519.5178,
  -63.89922,
  519.8635,
  -64.16969,
  97.78869,
  -296.2242,
  97.32874,
  -296.189,
  98.38185,
  -295.6939,
  98.15433,
  -296.0852,
  97.58721,
  -296.2755,
  97.45293,
  -296.4019,
  98.12043,
  -296.0403,
  97.63965,
  -296.1761,
  97.8474,
  -296.2304,
  97.23103,
  -296.4817,
  97.20521,
  -296.3142,
  96.66426,
  -296.4922,
  97.64149,
  -296.2845,
  97.561,
  -296.3621,
  96.79958,
  -296.5909,
  97.76905,
  -296.1624,
  98.05083,
  -295.9063,
  97.3813,
  -296.1327,
  97.12123,
  -296.1629,
  97.49383,
  -296.0043,
  97.76391,
  -295.54,
  97.47395,
  -295.7597,
  98.33752,
  -295.7967,
  97.64616,
  -296.1936,
  97.29415,
  -296.1773,
  97.52258,
  -296.2489,
  97.32834,
  -296.2009,
  97.53976,
  -295.9153,
  96.69438,
  -296.601,
  97.69356,
  -296.1923,
  97.36287,
  -296.2824,
  96.77269,
  -296.7282,
  97.28857,
  -296.4164,
  98.04126,
  -296.1071,
  97.46051,
  -296.3786,
  97.36913,
  -296.1954,
  98.26553,
  -295.5973,
  98.00439,
  -296.0436,
  97.85672,
  -296.1787,
  98.1736,
  -295.9427,
  98.2467,
  -295.9775,
  98.25191,
  -295.9647,
  97.86069,
  -296.1624,
  97.22234,
  -296.3065,
  96.79589,
  -296.4549,
  97.05755,
  -296.2964,
  97.75378,
  -296.1591,
  97.54385,
  -296.4293,
  96.72215,
  -296.6262,
  96.59352,
  -296.5553,
  97.89097,
  -295.6678,
  97.46032,
  -296.1545,
  96.95181,
  -296.4969,
  96.97573,
  -296.4148,
  98.31319,
  -295.7444,
  97.85769,
  -296.1917,
  97.29788,
  -296.3519,
  98.16043,
  -295.8747,
  97.71295,
  -295.9031,
  97.78703,
  -296.0421,
  97.70956,
  -296.1366,
  97.41636,
  -296.2334,
  97.15981,
  -296.4283,
  97.7081,
  -295.8509,
  97.59474,
  -296.1248,
  97.34794,
  -296.389,
  97.02536,
  -296.5974,
  97.05659,
  -296.5301,
  97.37784,
  -296.1984,
  97.18707,
  -296.4121,
  96.63385,
  -296.6116,
  97.01777,
  -296.5601,
  98.09141,
  -296.124,
  97.38354,
  -296.2957,
  96.76901,
  -296.6136,
  97.75146,
  -295.9933,
  98.05903,
  -295.8178,
  97.27544,
  -296.2375,
  97.05018,
  -296.4036,
  97.89421,
  -296.0703,
  98.05622,
  -295.8625,
  97.71998,
  -296.1046,
  97.31636,
  -296.2448,
  97.38177,
  -296.0984,
  98.11709,
  -295.781,
  97.91559,
  -295.9578,
  97.82832,
  -296.0008,
  96.89853,
  -296.3491,
  96.97137,
  -296.3645,
  97.74601,
  -296.1007,
  97.58506,
  -296.2989,
  97.36658,
  -296.3735,
  96.63857,
  -296.7162,
  97.21918,
  -296.3956,
  97.61425,
  -296.2461,
  97.08059,
  -296.4693,
  96.48267,
  -296.786,
  97.20245,
  -296.4005,
  97.75945,
  -295.9477,
  97.44152,
  -296.1701,
  96.75069,
  -296.5128,
  97.06865,
  -296.2719,
  97.93751,
  -295.7009,
  97.52421,
  -296.1108,
  97.05876,
  -296.3203,
  97.92332,
  -295.6617,
  98.29586,
  -295.5572,
  97.52566,
  -296.0786,
  97.03057,
  -296.3272,
  97.22793,
  -296.0028,
  98.0322,
  -295.481,
  97.80647,
  -295.6678,
  97.6408,
  -295.7863,
  97.24112,
  -296.3152,
  97.14822,
  -296.0674,
  97.95609,
  -295.8737,
  97.57742,
  -296.2065,
  97.1929,
  -296.5404,
  96.63118,
  -296.616,
  97.22211,
  -296.1705,
  97.52509,
  -295.9342,
  97.35456,
  -295.9013,
  96.46004,
  -296.5614,
  96.06716,
  -296.7097,
  97.10645,
  -296.1999,
  97.35378,
  -296.1528,
  97.02036,
  -296.4702,
  96.73281,
  -296.4454,
  97.7626,
  -295.9407,
  97.68365,
  -296.1871,
  97.16684,
  -296.35,
  96.58839,
  -296.5199,
  97.44777,
  -295.8601,
  97.89383,
  -295.9692,
  97.34893,
  -295.8603,
  96.77998,
  -296.4373,
  97.46515,
  -296.0812,
  98.02604,
  -295.855,
  97.63116,
  -296.0759,
  96.96819,
  -296.3794,
  97.7562,
  -295.9253,
  98.05122,
  -295.9433,
  97.88132,
  -296.0829,
  97.33701,
  -296.1543,
  98.09096,
  -295.7138,
  98.37474,
  -295.6791,
  97.80466,
  -295.8145,
  97.38881,
  -295.8855,
  96.94583,
  -296.2391,
  97.43784,
  -295.9374,
  97.92736,
  -295.7077,
  97.54253,
  -296.0428,
  97.15142,
  -296.2413,
  97.04242,
  -296.5592,
  97.51492,
  -296.1449,
  97.87137,
  -295.8214,
  97.12134,
  -296.1765,
  96.77264,
  -296.5127,
  96.27258,
  -296.8915,
  97.27122,
  -296.3507,
  97.25357,
  -296.1627,
  96.96644,
  -296.318,
  96.35323,
  -296.6678,
  97.34989,
  -296.1579,
  97.47594,
  -296.0561,
  97.17244,
  -296.2006,
  96.59775,
  -296.5071,
  97.71026,
  -296.0652,
  97.99982,
  -295.7615,
  97.31155,
  -296.0033,
  96.79822,
  -296.5331,
  97.69839,
  -295.8829,
  97.84579,
  -295.7346,
  97.47203,
  -296.0498,
  97.28355,
  -296.1713,
  98.36678,
  -295.7506,
  98.2817,
  -295.6772,
  97.89639,
  -295.9938,
  97.2075,
  -296.2619,
  97.29594,
  -296.3711,
  98.338,
  -295.7036,
  97.97358,
  -295.4991,
  97.22012,
  -295.9013,
  96.79734,
  -296.4706,
  97.73474,
  -296.0563,
  97.94424,
  -295.6853,
  97.50318,
  -295.9117,
  96.96052,
  -296.4188,
  97.00439,
  -296.3031,
  97.66106,
  -295.9341,
  97.8169,
  -295.8142,
  97.14977,
  -296.3469,
  96.90929,
  -296.411,
  97.10127,
  -296.2833,
  97.82673,
  -295.9328,
  97.45603,
  -295.9498,
  97.01398,
  -296.4095,
  96.70923,
  -296.361,
  97.00425,
  -296.3985,
  97.46593,
  -296.1134,
  96.9705,
  -296.1484,
  96.5014,
  -296.4117,
  96.67751,
  -296.5492,
  97.7601,
  -295.9779,
  97.27563,
  -296.305,
  96.83874,
  -296.4366,
  96.7336,
  -296.592,
  97.74578,
  -295.889,
  97.53532,
  -295.9297,
  96.83316,
  -296.2943,
  96.36259,
  -296.543,
  97.82459,
  -295.5595,
  97.66631,
  -295.6704,
  97.01443,
  -296.0492,
  96.88815,
  -296.3658,
  98.21601,
  -295.7728,
  97.84743,
  -295.8235,
  97.49265,
  -296.182,
  96.90064,
  -296.0414,
  97.88149,
  -295.6014,
  98.0454,
  -295.4908,
  97.43337,
  -295.5543,
  97.0279,
  -295.963,
  97.08794,
  -296.0395,
  98.05678,
  -295.8142,
  97.71618,
  -296.0334,
  97.22964,
  -295.9255,
  97.01805,
  -295.8551,
  97.19071,
  -295.6167,
  97.75681,
  -295.5001,
  97.47328,
  -295.9464,
  97.15999,
  -296.1302,
  97.35798,
  -296.4061,
  97.72429,
  -295.6256,
  97.24415,
  -295.8925,
  97.03094,
  -296.1269,
  96.86119,
  -296.2278,
  97.34718,
  -296.0101,
  97.32163,
  -296.0671,
  97.31638,
  -296.2912,
  96.91081,
  -296.2622,
  97.33044,
  -296.303,
  97.54316,
  -296.2542,
  97.53467,
  -296.1557,
  96.93607,
  -296.3135,
  96.45867,
  -296.2083,
  97.24282,
  -295.7905,
  97.45887,
  -295.6709,
  97.17267,
  -296.1236,
  96.7204,
  -296.5245,
  96.55636,
  -296.5439,
  97.4826,
  -295.7147,
  97.53072,
  -296.0448,
  96.83765,
  -296.1774,
  96.29567,
  -296.2517,
  97.70084,
  -295.9308,
  97.77848,
  -295.9388,
  97.18681,
  -296.107,
  96.91164,
  -296.3659,
  98.05626,
  -295.5709,
  97.94788,
  -295.6319,
  97.12635,
  -296.1338,
  96.92491,
  -296.517,
  97.48251,
  -296.073,
  97.98521,
  -295.615,
  97.4288,
  -295.7115,
  97.02055,
  -296.1152,
  97.78353,
  -295.864,
  98.02917,
  -295.9082,
  97.60637,
  -296.2098,
  97.39066,
  -296.0716,
  97.53774,
  -296.1299,
  98.32913,
  -295.7413,
  98.21963,
  -295.7722,
  97.7472,
  -296.0104,
  96.93062,
  -296.3942,
  98.11864,
  -295.8645,
  98.04227,
  -296.0215,
  97.29257,
  -296.2806,
  97.0612,
  -296.3119,
  97.13141,
  -296.4107,
  97.71686,
  -296.0036,
  97.88005,
  -296.0022,
  97.63915,
  -296.061,
  96.98928,
  -296.2577,
  97.16733,
  -296.2228,
  97.29404,
  -296.1646,
  97.3277,
  -296.0378,
  97.11646,
  -296.2477,
  96.80464,
  -296.2905,
  97.10436,
  -296.4114,
  97.58086,
  -296.1209,
  97.41631,
  -296.2105,
  96.98595,
  -296.3861,
  97.10445,
  -296.3289,
  97.6022,
  -296.1227,
  97.60061,
  -296.1835,
  97.05012,
  -296.4809,
  96.76064,
  -296.4977,
  97.83485,
  -296.0731,
  97.81599,
  -295.8578,
  97.35137,
  -296.3195,
  96.69047,
  -296.5394,
  97.58719,
  -296.1728,
  97.96935,
  -296.0722,
  97.67069,
  -296.2474,
  97.07877,
  -296.2807,
  97.93981,
  -295.828,
  98.20421,
  -295.8502,
  97.65548,
  -296.0493,
  97.12508,
  -296.4438,
  97.78471,
  -296.129,
  98.15974,
  -295.8127,
  97.89939,
  -296.0409,
  97.28072,
  -296.2708,
  97.14658,
  -296.1388,
  98.13809,
  -295.6744,
  98.02993,
  -295.956,
  -159.5753,
  -151.056,
  -159.8442,
  -150.7696,
  -158.8566,
  -151.3106,
  -159.3669,
  -151.4404,
  -159.5549,
  -151.0313,
  -159.8745,
  -150.8103,
  -159.2631,
  -151.3515,
  -159.6363,
  -151.0944,
  -159.5449,
  -151.1807,
  -160.1561,
  -150.8403,
  -159.7189,
  -150.6569,
  -160.3537,
  -150.4522,
  -159.6545,
  -151.1141,
  -159.896,
  -151.1002,
  -160.4542,
  -150.487,
  -159.4793,
  -151.1906,
  -159.2237,
  -151.452,
  -159.7668,
  -150.9466,
  -159.838,
  -150.917,
  -159.8699,
  -151.1027,
  -159.1809,
  -151.1505,
  -159.4951,
  -150.6344,
  -158.9461,
  -151.5694,
  -159.5208,
  -151.1863,
  -159.8704,
  -150.8813,
  -159.6548,
  -150.9726,
  -159.7053,
  -150.9369,
  -159.5497,
  -150.9323,
  -160.5407,
  -150.5939,
  -159.7245,
  -151.0362,
  -159.8737,
  -150.9288,
  -160.5305,
  -150.5098,
  -159.9261,
  -150.837,
  -159.3611,
  -151.3785,
  -159.901,
  -150.983,
  -159.8345,
  -150.7394,
  -158.8983,
  -151.4934,
  -159.2633,
  -151.2564,
  -159.4779,
  -151.1526,
  -159.2392,
  -151.3902,
  -159.1556,
  -151.4754,
  -159.1915,
  -151.5301,
  -159.6111,
  -151.1187,
  -159.9961,
  -150.776,
  -160.3463,
  -150.4342,
  -160.1295,
  -150.5781,
  -159.6156,
  -151.2132,
  -159.8691,
  -151.029,
  -160.4629,
  -150.373,
  -160.4611,
  -150.3869,
  -159.2289,
  -151.0305,
  -159.8365,
  -150.8581,
  -160.3438,
  -150.6961,
  -160.1952,
  -150.5247,
  -158.8988,
  -151.2358,
  -159.5175,
  -151.1865,
  -159.9324,
  -150.8677,
  -159.2141,
  -151.304,
  -159.5501,
  -151.0616,
  -159.3909,
  -151.1672,
  -159.528,
  -151.1436,
  -159.6626,
  -151.0444,
  -159.9324,
  -150.8669,
  -159.2946,
  -151.1143,
  -159.7832,
  -151.0156,
  -159.9223,
  -150.903,
  -160.2597,
  -150.7274,
  -160.1858,
  -150.7638,
  -159.6952,
  -150.9668,
  -160.0445,
  -150.8033,
  -160.4398,
  -150.3577,
  -160.1655,
  -150.5947,
  -159.2763,
  -151.2916,
  -159.9689,
  -150.8063,
  -160.4188,
  -150.5492,
  -159.5071,
  -151.0965,
  -159.1609,
  -151.2144,
  -159.7818,
  -150.7789,
  -160.1528,
  -150.5648,
  -159.4523,
  -151.12,
  -159.3009,
  -151.3186,
  -159.4922,
  -150.9993,
  -159.7693,
  -150.8343,
  -159.7784,
  -150.8495,
  -159.0826,
  -151.3677,
  -159.3484,
  -151.3546,
  -159.395,
  -151.0711,
  -160.0476,
  -150.6091,
  -160.16,
  -150.5794,
  -159.4367,
  -151.1955,
  -159.6927,
  -151.1132,
  -159.9281,
  -150.7815,
  -160.6092,
  -150.4747,
  -160.0469,
  -150.835,
  -159.7333,
  -151.0829,
  -160.1181,
  -150.79,
  -160.6676,
  -150.4061,
  -159.7859,
  -150.6564,
  -159.2971,
  -151.0398,
  -159.7015,
  -150.8214,
  -160.353,
  -150.458,
  -159.7424,
  -150.7662,
  -159.0559,
  -151.3986,
  -159.8252,
  -150.9308,
  -160.1383,
  -150.5707,
  -159.2727,
  -151.1882,
  -158.9387,
  -151.6275,
  -159.5693,
  -151.1931,
  -159.9871,
  -150.5307,
  -159.8051,
  -150.7315,
  -159.1679,
  -151.3155,
  -159.3691,
  -150.9165,
  -159.5189,
  -150.9754,
  -159.7981,
  -150.7984,
  -159.6397,
  -150.7018,
  -159.3668,
  -151.2442,
  -159.6511,
  -151.1514,
  -160.0332,
  -150.7334,
  -160.4106,
  -150.3605,
  -159.922,
  -150.8571,
  -159.5162,
  -151.0934,
  -159.5098,
  -150.7048,
  -160.4108,
  -150.1807,
  -160.6167,
  -150.0302,
  -159.8973,
  -150.6145,
  -159.6547,
  -150.9578,
  -160.1127,
  -150.8024,
  -160.3997,
  -150.5377,
  -159.3497,
  -151.0634,
  -159.4946,
  -151.0689,
  -160.0249,
  -150.8109,
  -160.4917,
  -150.2919,
  -159.3925,
  -150.9324,
  -159.4914,
  -151.2206,
  -160.0259,
  -150.7128,
  -160.3956,
  -150.4727,
  -159.6155,
  -151.0434,
  -158.8752,
  -151.3251,
  -159.6758,
  -151.1552,
  -160.0811,
  -150.6997,
  -159.376,
  -151.1622,
  -159.1531,
  -151.3924,
  -159.4625,
  -151.11,
  -159.7772,
  -150.8064,
  -158.7505,
  -151.4796,
  -158.949,
  -151.3332,
  -159.3333,
  -151.2978,
  -159.615,
  -150.9082,
  -160.2664,
  -150.5059,
  -159.6982,
  -150.9117,
  -158.8774,
  -151.366,
  -159.771,
  -151.0866,
  -160.1737,
  -150.8866,
  -160.4034,
  -150.7858,
  -159.7424,
  -150.9705,
  -159.4066,
  -151.232,
  -159.8545,
  -150.7832,
  -160.576,
  -150.5956,
  -160.7211,
  -150.2613,
  -159.8564,
  -150.8338,
  -159.9333,
  -150.6796,
  -160.1923,
  -150.6686,
  -160.7532,
  -150.2539,
  -159.5755,
  -150.8806,
  -159.6148,
  -151.0584,
  -159.9585,
  -150.7668,
  -160.5218,
  -150.4454,
  -159.4046,
  -151.1711,
  -159.3498,
  -151.3922,
  -159.7742,
  -150.867,
  -160.342,
  -150.4261,
  -159.6405,
  -151.113,
  -159.1746,
  -151.277,
  -159.5016,
  -150.8441,
  -160.0134,
  -150.7788,
  -158.9107,
  -151.4305,
  -159.0125,
  -151.3852,
  -159.4636,
  -151.3605,
  -159.7801,
  -150.8222,
  -159.7618,
  -150.847,
  -158.8661,
  -151.3208,
  -159.1015,
  -151.1644,
  -159.7196,
  -150.8836,
  -160.1387,
  -150.8561,
  -159.5336,
  -151.2124,
  -159.1216,
  -151.144,
  -159.8014,
  -150.8593,
  -160.004,
  -150.7519,
  -160.0239,
  -150.6107,
  -159.3469,
  -151.0133,
  -159.2461,
  -151.3151,
  -159.8407,
  -150.7392,
  -160.1952,
  -150.6904,
  -159.9751,
  -150.7831,
  -159.2807,
  -151.3264,
  -159.3651,
  -150.9247,
  -159.9358,
  -150.7891,
  -160.1823,
  -150.4528,
  -160.1283,
  -150.7121,
  -159.5903,
  -151.0083,
  -160.0689,
  -150.4069,
  -160.5502,
  -150.4467,
  -160.3696,
  -150.526,
  -159.435,
  -151.2276,
  -159.9808,
  -150.9123,
  -160.3083,
  -150.5617,
  -160.4296,
  -150.6441,
  -159.3893,
  -151.0542,
  -159.5983,
  -151.002,
  -160.0293,
  -150.5303,
  -160.2553,
  -150.1543,
  -158.8923,
  -151.1263,
  -159.1369,
  -151.091,
  -159.8124,
  -150.6378,
  -160.0755,
  -150.6192,
  -158.9347,
  -151.428,
  -159.3941,
  -151.2222,
  -159.6356,
  -150.8062,
  -159.7092,
  -150.4977,
  -158.8931,
  -151.2256,
  -159.1867,
  -151.3311,
  -159.4607,
  -150.8288,
  -160.064,
  -150.7285,
  -159.9402,
  -150.561,
  -159.1169,
  -151.44,
  -159.4025,
  -151.0716,
  -159.8232,
  -150.5743,
  -159.7997,
  -150.3129,
  -159.5323,
  -150.5271,
  -159.259,
  -150.9978,
  -159.6483,
  -150.8994,
  -160.1189,
  -150.8542,
  -159.9604,
  -150.9245,
  -159.1408,
  -151.2771,
  -159.4399,
  -150.8048,
  -160.0106,
  -150.7139,
  -160.069,
  -150.3994,
  -159.4946,
  -150.9972,
  -159.7118,
  -150.8352,
  -159.9066,
  -150.8299,
  -160.2222,
  -150.4391,
  -159.9428,
  -150.7251,
  -159.7618,
  -151.0687,
  -159.6164,
  -150.9538,
  -160.0081,
  -150.4258,
  -160.3234,
  -150.1297,
  -159.5866,
  -150.7717,
  -159.3314,
  -150.7453,
  -159.904,
  -150.7627,
  -160.3278,
  -150.4672,
  -160.4876,
  -150.2093,
  -159.5134,
  -150.755,
  -159.7134,
  -150.8428,
  -160.237,
  -150.4857,
  -160.5107,
  -150.0064,
  -159.4239,
  -151.0585,
  -159.3766,
  -151.1173,
  -159.8709,
  -150.7911,
  -160.1535,
  -150.5901,
  -158.974,
  -151.1843,
  -159.0911,
  -151.2588,
  -159.9265,
  -150.8304,
  -160.2613,
  -150.6348,
  -159.623,
  -151.0415,
  -159.1621,
  -151.1248,
  -159.5452,
  -151.0539,
  -159.8356,
  -150.6929,
  -159.4138,
  -151.1252,
  -159.1651,
  -151.3237,
  -159.6304,
  -150.9727,
  -159.7144,
  -150.9159,
  -159.6232,
  -150.9683,
  -159.0288,
  -151.3217,
  -158.998,
  -151.4302,
  -159.4501,
  -151.0131,
  -160.0647,
  -150.5987,
  -159.1423,
  -151.3393,
  -159.2105,
  -151.3637,
  -159.9233,
  -150.6507,
  -159.8112,
  -150.5595,
  -160.1331,
  -150.728,
  -159.5463,
  -150.9965,
  -159.2473,
  -151.1902,
  -159.6563,
  -150.9076,
  -160.1887,
  -150.6232,
  -159.9769,
  -150.624,
  -159.6635,
  -150.8266,
  -159.6779,
  -151.006,
  -160.1221,
  -150.6633,
  -160.399,
  -150.4584,
  -160.091,
  -150.6491,
  -159.6495,
  -151.1001,
  -159.8651,
  -151.0924,
  -160.0594,
  -150.7236,
  -160.0002,
  -150.7605,
  -159.5056,
  -151.0237,
  -159.5864,
  -151.0447,
  -160.1853,
  -150.7485,
  -160.277,
  -150.4682,
  -159.565,
  -151.2099,
  -159.4134,
  -151.1357,
  -159.9271,
  -150.9354,
  -160.3671,
  -150.4943,
  -159.596,
  -150.9446,
  -159.3126,
  -151.2952,
  -159.7871,
  -150.9179,
  -159.986,
  -150.584,
  -159.2834,
  -151.0526,
  -159.0497,
  -151.5026,
  -159.472,
  -151.0029,
  -160.0851,
  -150.7533,
  -159.437,
  -151.271,
  -159.0852,
  -151.5798,
  -159.5884,
  -151.2727,
  -159.7547,
  -150.8745,
  -159.5541,
  -150.6815,
  -158.8684,
  -151.309,
  -159.2301,
  -151.3931,
  -156.3122,
  60.97182,
  -156.2296,
  61.60086,
  -156.204,
  60.21061,
  -156.317,
  60.64019,
  -156.1541,
  61.12182,
  -156.2485,
  61.38223,
  -156.2775,
  60.68825,
  -156.2997,
  61.08392,
  -156.4626,
  60.82326,
  -156.2463,
  61.5943,
  -155.9413,
  61.43772,
  -156.123,
  62.10432,
  -156.3216,
  61.10249,
  -156.396,
  61.25625,
  -156.2361,
  62.01009,
  -156.2448,
  60.8589,
  -156.3278,
  60.64494,
  -156.1657,
  61.3422,
  -155.9646,
  61.44635,
  -156.0641,
  61.0776,
  -155.7801,
  60.72212,
  -156.1137,
  61.14292,
  -156.2556,
  60.31506,
  -156.3004,
  60.95322,
  -156.2388,
  61.56037,
  -156.638,
  61.50607,
  -156.1777,
  61.6045,
  -156.2229,
  61.18901,
  -156.0494,
  61.84082,
  -156.3438,
  60.88774,
  -156.2688,
  61.55966,
  -156.1281,
  62.09147,
  -156.1815,
  61.44614,
  -156.4368,
  60.63417,
  -156.3748,
  61.33541,
  -156.1995,
  61.3068,
  -156.2738,
  60.18823,
  -156.2747,
  60.80523,
  -156.455,
  60.97504,
  -156.418,
  60.57426,
  -156.3904,
  60.48987,
  -156.4926,
  60.42589,
  -156.4752,
  60.86536,
  -156.0824,
  61.41297,
  -156.1433,
  61.895,
  -156.1274,
  61.62483,
  -156.3523,
  61.04505,
  -156.3379,
  61.32596,
  -156.1109,
  62.05192,
  -156.127,
  62.11165,
  -156.2081,
  60.72221,
  -156.2256,
  61.10239,
  -156.0993,
  61.79805,
  -156.3651,
  61.65931,
  -156.4466,
  60.40869,
  -156.4286,
  60.76149,
  -156.271,
  61.45647,
  -156.3233,
  60.64961,
  -156.3336,
  60.85413,
  -156.3981,
  60.83621,
  -156.3652,
  60.85213,
  -156.4741,
  61.13188,
  -156.2386,
  61.46095,
  -156.3449,
  60.80409,
  -156.2088,
  61.03249,
  -156.2039,
  61.43161,
  -156.279,
  61.85101,
  -156.2075,
  61.70988,
  -156.2173,
  61.38007,
  -156.1769,
  61.56014,
  -156.2914,
  62.26931,
  -156.2645,
  61.71023,
  -156.4683,
  60.76343,
  -156.2199,
  61.35083,
  -156.138,
  62.14041,
  -156.1281,
  60.94948,
  -156.2972,
  60.59846,
  -156.2643,
  61.14961,
  -156.3033,
  61.76156,
  -156.3022,
  60.82872,
  -156.2173,
  60.635,
  -156.3181,
  60.96868,
  -156.264,
  61.37223,
  -156.2745,
  61.12509,
  -156.3638,
  60.57541,
  -156.534,
  60.87111,
  -156.3183,
  60.85168,
  -156.1627,
  61.60418,
  -156.1301,
  61.76431,
  -156.3049,
  60.95821,
  -156.4053,
  61.19631,
  -156.6694,
  61.32633,
  -156.2725,
  62.23458,
  -156.2569,
  61.60439,
  -156.3606,
  61.18218,
  -156.2821,
  61.69334,
  -156.2231,
  62.31902,
  -156.0915,
  61.70776,
  -156.2842,
  60.82582,
  -156.4126,
  61.22937,
  -156.2322,
  61.92372,
  -155.9951,
  61.60791,
  -156.3463,
  60.69013,
  -156.4769,
  61.29008,
  -156.2659,
  61.87918,
  -156.2869,
  60.68668,
  -156.3794,
  60.44969,
  -156.2115,
  61.22919,
  -156.2639,
  61.68506,
  -156.0367,
  61.46889,
  -156.088,
  60.69756,
  -156.1989,
  60.93823,
  -156.0862,
  61.29526,
  -156.1468,
  61.52274,
  -156.1495,
  61.62093,
  -156.5563,
  60.65094,
  -156.4932,
  61.10424,
  -156.2184,
  61.89665,
  -156.2005,
  62.30777,
  -156.0207,
  61.40055,
  -156.2782,
  61.11736,
  -156.5152,
  61.26314,
  -156.3163,
  61.96194,
  -155.9395,
  62.38012,
  -156.0824,
  61.47819,
  -156.2175,
  61.37957,
  -156.1799,
  61.8296,
  -156.1254,
  62.03448,
  -156.2332,
  60.87391,
  -156.4449,
  61.05061,
  -156.3611,
  61.58053,
  -156.0133,
  62.29456,
  -156.1131,
  60.97142,
  -156.3442,
  60.85786,
  -156.2159,
  61.36815,
  -156.121,
  61.98035,
  -156.1904,
  61.12873,
  -156.3377,
  60.44817,
  -156.1447,
  61.05581,
  -156.1639,
  61.71321,
  -156.1713,
  60.85197,
  -156.346,
  60.56237,
  -156.3757,
  61.00425,
  -156.2418,
  61.37833,
  -156.2677,
  60.5645,
  -156.4814,
  60.38969,
  -156.3914,
  60.92184,
  -156.1887,
  61.35447,
  -156.2352,
  61.92103,
  -156.2355,
  61.1375,
  -156.4091,
  60.65068,
  -156.3253,
  61.37467,
  -156.0203,
  61.55311,
  -156.2401,
  61.66151,
  -156.2541,
  61.16217,
  -156.1755,
  60.79037,
  -156.2399,
  61.619,
  -156.1552,
  62.19656,
  -156.0897,
  62.48482,
  -156.4166,
  61.40149,
  -156.2775,
  61.32256,
  -156.109,
  61.93466,
  -156.2122,
  62.47007,
  -156.2192,
  61.43716,
  -156.2824,
  61.07066,
  -156.2692,
  61.62128,
  -156.1115,
  62.03065,
  -156.3342,
  61.06398,
  -156.4615,
  60.64377,
  -156.1465,
  61.51046,
  -156.3663,
  61.93159,
  -156.2309,
  60.75467,
  -156.2435,
  60.64568,
  -156.3887,
  61.19595,
  -156.2997,
  61.49468,
  -156.3319,
  60.3014,
  -156.2673,
  60.32854,
  -156.2816,
  60.90058,
  -156.2039,
  61.47077,
  -156.151,
  61.41646,
  -156.2354,
  60.09729,
  -156.3259,
  60.58216,
  -156.3019,
  61.33139,
  -156.1944,
  61.6343,
  -156.2817,
  60.83073,
  -156.3018,
  60.65822,
  -156.2444,
  61.29596,
  -156.283,
  61.81829,
  -156.2085,
  61.75756,
  -156.1054,
  61.11059,
  -156.2883,
  60.73642,
  -156.4905,
  61.21696,
  -156.22,
  61.79875,
  -156.1825,
  61.60145,
  -156.3149,
  60.96485,
  -156.2671,
  61.28434,
  -156.4542,
  61.62881,
  -155.9699,
  61.753,
  -156.1965,
  61.80108,
  -156.4046,
  61.00114,
  -156.2366,
  61.48104,
  -156.1427,
  62.12364,
  -156.3666,
  62.11037,
  -156.3599,
  60.9002,
  -156.3271,
  61.4615,
  -156.2895,
  61.93434,
  -156.1853,
  62.18913,
  -156.1513,
  60.84865,
  -156.2799,
  60.9063,
  -156.4671,
  61.85273,
  -156.1578,
  62.27953,
  -156.1683,
  60.85818,
  -156.14,
  60.989,
  -156.1002,
  61.66505,
  -156.0911,
  61.98956,
  -156.41,
  60.21362,
  -156.3469,
  60.7298,
  -156.508,
  61.27251,
  -156.0245,
  61.85633,
  -155.9647,
  60.61372,
  -156.0542,
  60.45575,
  -156.0313,
  60.72956,
  -156.1626,
  61.43996,
  -156.267,
  61.38025,
  -156.304,
  60.41305,
  -156.5337,
  60.81052,
  -156.1409,
  61.42868,
  -156.1771,
  61.80222,
  -155.8043,
  61.31782,
  -155.9919,
  60.86089,
  -156.2068,
  61.10007,
  -156.3362,
  61.75541,
  -156.1693,
  61.42267,
  -156.2035,
  60.70033,
  -156.0928,
  61.21303,
  -156.2142,
  61.37637,
  -156.0755,
  61.43955,
  -156.4524,
  61.32595,
  -156.4838,
  61.25901,
  -156.2845,
  61.52032,
  -156.0466,
  61.83622,
  -156.1601,
  61.30779,
  -156.3762,
  61.15352,
  -156.426,
  61.1028,
  -156.3849,
  61.59282,
  -155.9084,
  62.59351,
  -156.0287,
  61.56754,
  -156.1687,
  60.88136,
  -156.0026,
  61.52438,
  -156.1835,
  62.02795,
  -156.3012,
  62.25141,
  -156.265,
  60.9658,
  -156.3559,
  61.15923,
  -155.8962,
  61.70184,
  -155.9637,
  62.32875,
  -156.1478,
  60.94257,
  -156.2222,
  60.89307,
  -156.0937,
  61.4575,
  -156.0565,
  61.88727,
  -155.9588,
  60.42134,
  -156.1157,
  60.64515,
  -156.2126,
  61.34368,
  -156.3899,
  61.904,
  -156.3452,
  61.15543,
  -156.3162,
  60.64511,
  -156.085,
  61.00838,
  -156.1968,
  61.37259,
  -156.3166,
  61.01377,
  -156.325,
  60.59057,
  -156.311,
  61.19287,
  -156.1496,
  61.25079,
  -156.2888,
  61.13423,
  -156.2615,
  60.40107,
  -156.3503,
  60.61295,
  -156.2354,
  61.12474,
  -156.1422,
  61.75652,
  -156.1655,
  60.63294,
  -156.3454,
  60.55783,
  -156.2739,
  61.55257,
  -156.0377,
  61.70259,
  -156.2817,
  61.6818,
  -156.1323,
  61.01136,
  -156.2587,
  60.82043,
  -156.12,
  61.28264,
  -156.2292,
  61.75887,
  -156.1811,
  61.60903,
  -156.17,
  61.4217,
  -156.3202,
  61.20267,
  -156.2959,
  61.69818,
  -156.0684,
  62.03218,
  -156.2987,
  61.71641,
  -156.3264,
  61.16364,
  -156.3156,
  61.2961,
  -156.1386,
  61.69964,
  -156.1912,
  61.66279,
  -156.1746,
  61.07747,
  -156.2192,
  61.15613,
  -156.3277,
  61.73688,
  -156.2392,
  62.16626,
  -156.2009,
  61.0395,
  -156.2831,
  60.89991,
  -156.2838,
  61.47189,
  -156.1942,
  62.10273,
  -156.1962,
  61.08724,
  -156.322,
  60.67172,
  -156.4576,
  61.22912,
  -156.1799,
  61.78299,
  -156.1095,
  60.61647,
  -156.347,
  60.44319,
  -156.1804,
  61.04473,
  -156.2036,
  61.60485,
  -156.2803,
  60.91468,
  -156.2766,
  60.46131,
  -156.3233,
  60.86908,
  -156.4309,
  61.38142,
  -156.2627,
  61.35357,
  -156.1932,
  60.41601,
  -156.3184,
  60.76946,
  -9.135457,
  133.9586,
  -8.805316,
  134.0869,
  -9.868482,
  133.6278,
  -9.489536,
  133.8985,
  -8.987088,
  134.0178,
  -8.723711,
  134.1036,
  -9.53311,
  133.7651,
  -9.119905,
  134.0729,
  -9.249376,
  134.0144,
  -8.629782,
  134.2586,
  -8.746415,
  134.2146,
  -8.151993,
  134.3008,
  -9.120995,
  133.9065,
  -8.922902,
  134.1882,
  -8.187552,
  134.3051,
  -9.226713,
  133.7906,
  -9.532727,
  133.846,
  -8.831526,
  134.0662,
  -8.688764,
  134.0803,
  -8.897079,
  134.0356,
  -9.106925,
  133.5064,
  -8.881607,
  133.7197,
  -9.799979,
  133.4803,
  -9.430359,
  133.9336,
  -8.81442,
  134.0843,
  -9.136968,
  133.8725,
  -9.019121,
  134.0368,
  -8.989437,
  134.0301,
  -8.125579,
  134.2711,
  -9.31231,
  133.6934,
  -8.806966,
  134.0987,
  -8.16414,
  134.3985,
  -8.764901,
  134.0555,
  -9.420671,
  133.9322,
  -8.914673,
  134.0726,
  -8.80621,
  133.9488,
  -9.966488,
  133.5118,
  -9.423043,
  133.9164,
  -9.296165,
  134.0191,
  -9.609938,
  133.7022,
  -9.57583,
  133.6908,
  -9.719948,
  133.782,
  -9.242886,
  133.8711,
  -8.692471,
  134.153,
  -8.183899,
  134.3146,
  -8.592274,
  134.0943,
  -9.220564,
  133.9922,
  -8.919509,
  134.1958,
  -8.304423,
  134.3871,
  -8.048967,
  134.2889,
  -9.350272,
  133.7011,
  -9.119423,
  134.1027,
  -8.604239,
  134.327,
  -8.476886,
  134.1008,
  -9.737669,
  133.7802,
  -9.289804,
  134.0424,
  -8.674558,
  134.1097,
  -9.509874,
  133.7612,
  -9.287728,
  133.9099,
  -9.344876,
  133.8847,
  -9.188583,
  133.9424,
  -8.980599,
  134.0559,
  -8.621697,
  134.0865,
  -9.239202,
  133.718,
  -9.108131,
  134.106,
  -8.747596,
  134.0628,
  -8.423133,
  134.3206,
  -8.525249,
  134.2829,
  -8.794627,
  133.8771,
  -8.538258,
  134.2548,
  -7.94551,
  134.3924,
  -8.3967,
  134.118,
  -9.382429,
  133.8927,
  -8.805926,
  134.1851,
  -8.32414,
  134.3753,
  -9.237949,
  133.8132,
  -9.493939,
  133.7967,
  -8.96174,
  134.1397,
  -8.517042,
  134.202,
  -9.320601,
  133.8153,
  -9.520817,
  133.7101,
  -9.145827,
  134.0511,
  -8.707321,
  134.1405,
  -8.703221,
  133.9795,
  -9.565619,
  133.6192,
  -9.395402,
  133.8661,
  -9.297282,
  133.9849,
  -8.531776,
  134.1879,
  -8.415919,
  134.1359,
  -9.183751,
  133.9201,
  -9.068003,
  134.0555,
  -8.93585,
  134.2405,
  -8.149835,
  134.3895,
  -8.640676,
  134.1178,
  -9.015725,
  134.0403,
  -8.537457,
  134.1986,
  -7.922197,
  134.4862,
  -8.683231,
  134.0953,
  -9.250403,
  133.8663,
  -8.841889,
  134.259,
  -8.248546,
  134.357,
  -8.671762,
  134.0713,
  -9.638009,
  133.7552,
  -9.117782,
  134.1291,
  -8.411471,
  134.2338,
  -9.192921,
  133.8328,
  -9.622111,
  133.4262,
  -9.139234,
  133.8022,
  -8.655613,
  134.1857,
  -8.745235,
  134.0441,
  -9.439394,
  133.5657,
  -9.028032,
  133.7777,
  -9.009732,
  133.9739,
  -8.56612,
  134.3319,
  -8.729308,
  134.0637,
  -9.545493,
  133.7805,
  -9.050832,
  134.0832,
  -8.492682,
  134.1663,
  -8.019179,
  134.3495,
  -8.774204,
  134.0196,
  -9.231211,
  134.0382,
  -8.774663,
  134.0178,
  -8.239791,
  134.4015,
  -7.688596,
  134.5113,
  -8.584228,
  134.1628,
  -8.707961,
  134.1896,
  -8.36748,
  134.3663,
  -8.13982,
  134.3588,
  -9.253383,
  133.7684,
  -9.136901,
  133.953,
  -8.618269,
  134.2423,
  -8.036895,
  134.3363,
  -9.10666,
  133.8333,
  -9.434401,
  133.8918,
  -8.748071,
  134.0543,
  -8.169525,
  134.2176,
  -9.04096,
  133.8567,
  -9.500818,
  133.7192,
  -8.914635,
  134.0752,
  -8.446165,
  134.2067,
  -9.217649,
  133.7216,
  -9.604208,
  133.706,
  -9.213058,
  133.9634,
  -8.750359,
  134.0827,
  -9.624093,
  133.4111,
  -9.703143,
  133.5078,
  -9.290584,
  133.8951,
  -9.043874,
  134.0296,
  -8.434718,
  134.2433,
  -9.06848,
  133.8798,
  -9.43577,
  133.8673,
  -8.964247,
  134.0642,
  -8.725204,
  134.2351,
  -8.422403,
  134.285,
  -9.001907,
  134.0414,
  -9.360645,
  133.8673,
  -8.78661,
  134.223,
  -8.145827,
  134.4519,
  -7.854006,
  134.621,
  -8.880251,
  134.2251,
  -8.749851,
  134.2243,
  -8.379904,
  134.4341,
  -8.007271,
  134.4532,
  -8.75352,
  133.9758,
  -9.063841,
  134.0796,
  -8.699822,
  134.2651,
  -8.030319,
  134.5267,
  -9.119692,
  133.9533,
  -9.381047,
  133.9124,
  -8.660367,
  134.1346,
  -8.229873,
  134.3952,
  -9.079798,
  133.6186,
  -9.480832,
  133.7843,
  -9.15014,
  133.908,
  -8.851923,
  134.181,
  -9.822231,
  133.6669,
  -9.80636,
  133.6657,
  -9.290484,
  133.9888,
  -8.652536,
  134.2036,
  -8.849488,
  134.0677,
  -9.98547,
  133.6276,
  -9.586432,
  133.7449,
  -8.944204,
  134.0852,
  -8.589804,
  134.2414,
  -9.38482,
  133.8985,
  -9.58559,
  133.6772,
  -8.98273,
  134.0061,
  -8.62752,
  134.3836,
  -8.60228,
  134.1926,
  -9.204787,
  133.938,
  -9.433572,
  133.7772,
  -8.881431,
  134.2329,
  -8.421125,
  134.1541,
  -8.618167,
  134.0373,
  -9.319454,
  133.9572,
  -8.813386,
  134.0133,
  -8.61704,
  134.3141,
  -8.395185,
  134.1332,
  -8.524384,
  134.2043,
  -9.170566,
  134.0323,
  -8.494421,
  134.069,
  -8.029476,
  134.4852,
  -8.134211,
  134.4672,
  -9.234982,
  133.8789,
  -8.89842,
  134.1585,
  -8.421836,
  134.3355,
  -8.168087,
  134.3884,
  -9.271252,
  133.7272,
  -9.333386,
  134.068,
  -8.664001,
  134.4273,
  -8.31499,
  134.3351,
  -9.475629,
  133.6161,
  -9.310398,
  133.7096,
  -8.687313,
  134.1859,
  -8.403937,
  134.2155,
  -9.86432,
  133.495,
  -9.538321,
  133.7955,
  -8.953585,
  134.0355,
  -8.446996,
  133.8113,
  -9.52275,
  133.6306,
  -9.63502,
  133.5925,
  -9.348933,
  134.1577,
  -8.730947,
  134.2247,
  -8.669488,
  134.1016,
  -9.704088,
  133.7331,
  -9.410659,
  133.9537,
  -8.623412,
  134.2572,
  -8.444605,
  134.1271,
  -8.811094,
  133.763,
  -9.162573,
  133.7394,
  -8.961413,
  134.1673,
  -8.749318,
  134.1645,
  -8.719611,
  134.0016,
  -9.341789,
  133.4451,
  -8.602629,
  133.9833,
  -8.647351,
  134.0918,
  -8.632836,
  134.1416,
  -8.772613,
  133.9892,
  -8.884159,
  133.9324,
  -8.787015,
  134.0805,
  -8.26565,
  134.2715,
  -8.722037,
  134.1129,
  -9.033588,
  134.0336,
  -9.081685,
  134.1096,
  -8.587768,
  134.3165,
  -7.905381,
  134.356,
  -8.792418,
  134.0167,
  -9.213684,
  133.8614,
  -8.688154,
  134.0137,
  -8.170286,
  134.3549,
  -8.135158,
  134.3636,
  -9.013107,
  133.6998,
  -9.085229,
  134.0964,
  -8.516309,
  134.2346,
  -7.908556,
  134.3448,
  -9.196762,
  133.8674,
  -9.229192,
  133.9246,
  -8.657224,
  134,
  -8.331236,
  134.1113,
  -9.51639,
  133.5718,
  -9.4511,
  133.6728,
  -8.732771,
  134.2286,
  -8.327967,
  134.4118,
  -8.923436,
  134.0251,
  -9.329226,
  133.7502,
  -9.028307,
  133.7716,
  -8.651619,
  134.1431,
  -9.165346,
  133.8029,
  -9.500083,
  133.8171,
  -9.119481,
  133.919,
  -8.74646,
  133.9271,
  -8.971452,
  133.9798,
  -9.642523,
  133.6467,
  -9.589424,
  133.7241,
  -9.173183,
  133.8998,
  -8.535812,
  134.2532,
  -9.504222,
  133.7561,
  -9.586291,
  133.8208,
  -8.488228,
  134.222,
  -8.580844,
  134.0997,
  -8.590674,
  134.2617,
  -9.141512,
  133.8366,
  -9.356075,
  133.7722,
  -8.876314,
  134.0787,
  -8.407894,
  134.2198,
  -8.556447,
  134.182,
  -8.768678,
  134.1294,
  -8.829388,
  134.1365,
  -8.569503,
  134.1093,
  -8.234684,
  134.1499,
  -8.549394,
  134.2115,
  -9.016842,
  133.9851,
  -8.93368,
  134.0353,
  -8.564446,
  134.1878,
  -8.619871,
  134.1311,
  -9.153317,
  133.8945,
  -9.270854,
  134.0921,
  -8.567855,
  134.2359,
  -8.251354,
  134.3268,
  -9.296835,
  133.9954,
  -9.218262,
  133.8025,
  -8.737812,
  134.2041,
  -8.178126,
  134.3913,
  -9.071939,
  133.7959,
  -9.529107,
  133.7968,
  -8.988797,
  134.1348,
  -8.477416,
  134.184,
  -9.30624,
  133.6021,
  -9.641342,
  133.7528,
  -9.181249,
  133.9558,
  -8.547865,
  134.1965,
  -9.269751,
  133.9094,
  -9.673532,
  133.6676,
  -9.368781,
  133.9689,
  -8.836574,
  134.1464,
  -8.701526,
  134.1147,
  -9.659003,
  133.5422,
  -9.477873,
  133.8292,
  96.64702,
  53.87895,
  96.86759,
  53.49522,
  95.89323,
  54.24051,
  96.33448,
  54.07492,
  96.62151,
  53.81536,
  96.89398,
  53.61079,
  96.24081,
  54.03342,
  96.68494,
  53.74918,
  96.5957,
  53.95713,
  97.04021,
  53.5111,
  96.77229,
  53.5672,
  97.37828,
  53.17188,
  96.64265,
  53.73263,
  96.94239,
  53.7731,
  97.38539,
  53.15443,
  96.40351,
  53.77769,
  96.25876,
  54.09082,
  96.80212,
  53.66111,
  96.89024,
  53.61305,
  96.68158,
  53.67017,
  96.39964,
  53.66671,
  96.56874,
  53.63207,
  95.85379,
  54.24902,
  96.50029,
  53.94798,
  96.97716,
  53.65685,
  96.64461,
  53.65199,
  96.73436,
  53.66461,
  96.67326,
  53.77733,
  97.47145,
  53.05394,
  96.40496,
  53.78531,
  96.93838,
  53.57451,
  97.43801,
  53.12495,
  96.86504,
  53.48197,
  96.41129,
  54.09932,
  96.97918,
  53.71471,
  96.82043,
  53.53782,
  95.90616,
  54.21993,
  96.29984,
  54.02094,
  96.64525,
  53.96315,
  96.17373,
  54.10739,
  96.10209,
  54.18088,
  96.13503,
  54.31259,
  96.61012,
  53.91549,
  96.96096,
  53.48646,
  97.31561,
  53.29549,
  96.94523,
  53.39967,
  96.52754,
  53.79864,
  96.84631,
  53.71458,
  97.40519,
  53.14158,
  97.46025,
  53.02666,
  96.29221,
  53.92485,
  96.78786,
  53.74121,
  97.19317,
  53.39726,
  96.9986,
  53.27936,
  96.0433,
  54.22172,
  96.58417,
  54.00617,
  96.98634,
  53.46666,
  96.18569,
  54.04127,
  96.52941,
  54.01624,
  96.3892,
  53.95347,
  96.46783,
  53.94199,
  96.76102,
  53.7792,
  96.9633,
  53.53269,
  96.42342,
  53.83627,
  96.81702,
  53.87919,
  96.92994,
  53.55653,
  97.22815,
  53.33337,
  97.16255,
  53.41538,
  96.76286,
  53.56822,
  97.0338,
  53.44678,
  97.46325,
  53.00691,
  97.04155,
  53.32346,
  96.35104,
  54.06827,
  96.8895,
  53.55029,
  97.3614,
  53.1877,
  96.44482,
  53.87259,
  96.24481,
  54.16481,
  96.74383,
  53.70443,
  97.14436,
  53.38289,
  96.38004,
  53.88499,
  96.12524,
  54.04486,
  96.62965,
  53.87481,
  97.06286,
  53.51779,
  96.73282,
  53.6448,
  96.1634,
  54.06758,
  96.52522,
  54.10102,
  96.46204,
  53.95407,
  97.00536,
  53.27327,
  97.11042,
  53.20876,
  96.49603,
  53.82591,
  96.71442,
  53.75773,
  96.94669,
  53.66817,
  97.53753,
  53.16065,
  96.9827,
  53.47435,
  96.73061,
  53.84836,
  97.15321,
  53.44464,
  97.61956,
  53.07003,
  96.90255,
  53.39827,
  96.42461,
  53.867,
  96.89398,
  53.6498,
  97.37128,
  53.23698,
  96.79183,
  53.54873,
  96.18315,
  54.25331,
  96.86581,
  53.90277,
  97.20206,
  53.30682,
  96.2476,
  53.90206,
  95.86059,
  54.09067,
  96.46753,
  53.77734,
  97.02757,
  53.5422,
  96.8905,
  53.67448,
  96.17626,
  53.98367,
  96.35218,
  53.96997,
  96.92174,
  53.79911,
  97.00765,
  53.49791,
  96.76988,
  53.53966,
  96.20673,
  54.10315,
  96.68922,
  53.87238,
  97.11374,
  53.4243,
  97.49072,
  53.15843,
  96.73139,
  53.54971,
  96.47629,
  54.00195,
  96.79929,
  53.60886,
  97.42571,
  53.07729,
  97.61314,
  52.92944,
  97.00909,
  53.4777,
  96.85353,
  53.6856,
  97.24443,
  53.31521,
  97.38966,
  53.24944,
  96.34148,
  53.79144,
  96.52309,
  53.89057,
  97.0727,
  53.54334,
  97.48786,
  53.03484,
  96.34961,
  53.72533,
  96.35938,
  54.04153,
  96.68723,
  53.48436,
  97.25336,
  53.18615,
  96.51708,
  53.67507,
  96.21527,
  54.06978,
  96.7085,
  53.62507,
  97.14545,
  53.29823,
  96.45296,
  53.76919,
  96.13883,
  54.08789,
  96.57083,
  53.81747,
  96.94221,
  53.54913,
  96.13799,
  54.07966,
  95.91902,
  54.21062,
  96.41119,
  53.9468,
  96.78959,
  53.69254,
  97.20551,
  53.45646,
  96.54154,
  53.6801,
  96.36398,
  54.09034,
  96.79597,
  53.75066,
  97.03465,
  53.5748,
  97.2161,
  53.38077,
  96.67397,
  53.69977,
  96.41595,
  54.03843,
  97.00555,
  53.62552,
  97.45506,
  53.2143,
  97.80662,
  52.9592,
  96.88012,
  53.70704,
  96.86877,
  53.68002,
  97.37357,
  53.37928,
  97.60499,
  53.05499,
  96.72742,
  53.64057,
  96.59653,
  54.00798,
  97.02154,
  53.53953,
  97.42753,
  53.08992,
  96.55828,
  53.88212,
  96.36878,
  54.03875,
  96.90504,
  53.56651,
  97.30447,
  53.25599,
  96.48523,
  53.65827,
  96.17878,
  54.04278,
  96.68509,
  53.75077,
  96.822,
  53.58644,
  95.97007,
  54.20083,
  95.95235,
  54.27504,
  96.52716,
  54.03114,
  96.92245,
  53.56248,
  96.82761,
  53.57005,
  95.96375,
  54.34246,
  96.3055,
  54.10231,
  96.79205,
  53.65866,
  97.07183,
  53.46865,
  96.46325,
  53.9838,
  96.23161,
  54.01941,
  96.80875,
  53.70501,
  97.12026,
  53.37077,
  97.15701,
  53.33998,
  96.57227,
  53.82545,
  96.3409,
  53.96688,
  96.90331,
  53.5849,
  97.17285,
  53.35528,
  96.98007,
  53.35673,
  96.52791,
  54.00579,
  96.81792,
  53.72931,
  97.1073,
  53.50181,
  97.20132,
  53.34257,
  97.07552,
  53.34497,
  96.70374,
  53.74261,
  97.06309,
  53.36117,
  97.46898,
  53.08167,
  97.55083,
  53.12767,
  96.53133,
  53.89431,
  96.95039,
  53.67654,
  97.2975,
  53.31109,
  97.39589,
  53.15074,
  96.37026,
  53.83324,
  96.76374,
  53.85136,
  97.19781,
  53.47216,
  97.38287,
  53.01285,
  96.13593,
  53.87077,
  96.42819,
  54.01876,
  96.8403,
  53.59753,
  97.14975,
  53.26606,
  95.85133,
  54.272,
  96.28233,
  54.01039,
  96.76755,
  53.66652,
  97.09746,
  53.00725,
  96.06603,
  53.86991,
  96.10011,
  53.95955,
  96.56047,
  54.00035,
  96.97103,
  53.4963,
  96.92615,
  53.44019,
  96.08788,
  54.20059,
  96.55474,
  54.00429,
  96.87663,
  53.56397,
  96.91508,
  53.49185,
  96.69376,
  53.698,
  96.40902,
  53.91849,
  96.69714,
  53.76483,
  96.9705,
  53.55806,
  96.88783,
  53.5592,
  96.18266,
  53.81021,
  96.71789,
  53.59085,
  97.03117,
  53.46511,
  97.02351,
  53.4139,
  96.68382,
  53.48247,
  96.57716,
  53.58493,
  96.82219,
  53.59773,
  97.21136,
  53.25978,
  96.86754,
  53.55514,
  96.73705,
  53.76072,
  96.72008,
  53.81272,
  97.18199,
  53.54074,
  97.57582,
  53.03568,
  96.68771,
  53.43079,
  96.55422,
  53.7734,
  96.94307,
  53.48628,
  97.52943,
  53.18549,
  97.47403,
  53.23972,
  96.47316,
  53.72628,
  96.75262,
  53.79195,
  97.16876,
  53.29689,
  97.64797,
  52.91267,
  96.43231,
  53.81736,
  96.58899,
  53.90601,
  96.91089,
  53.41924,
  97.18123,
  53.21349,
  96.01588,
  53.84572,
  96.18841,
  53.98294,
  96.9398,
  53.56201,
  97.41837,
  53.3959,
  96.73146,
  53.77011,
  96.19893,
  54.05309,
  96.51569,
  53.70632,
  96.80228,
  53.51662,
  96.42987,
  53.71776,
  96.18985,
  54.02875,
  96.58229,
  53.82766,
  96.76733,
  53.59195,
  96.64936,
  53.71112,
  95.96453,
  54.10201,
  96.19262,
  54.06142,
  96.68972,
  53.83073,
  97.08865,
  53.41349,
  96.21506,
  54.04187,
  96.21871,
  54.09161,
  97.00854,
  53.35272,
  97.01295,
  53.34519,
  97.14678,
  53.41835,
  96.49732,
  53.69056,
  96.43167,
  53.97525,
  96.91331,
  53.62441,
  97.18999,
  53.36354,
  96.9203,
  53.4687,
  96.77972,
  53.54855,
  96.87666,
  53.59909,
  97.11201,
  53.4137,
  97.3637,
  53.1273,
  97.10474,
  53.41452,
  96.64366,
  53.7933,
  96.89482,
  53.71804,
  97.16553,
  53.38324,
  96.99638,
  53.44564,
  96.56923,
  53.69914,
  96.70252,
  53.97455,
  97.19132,
  53.4897,
  97.35705,
  53.13908,
  96.51,
  53.87242,
  96.49865,
  53.88786,
  96.92491,
  53.57679,
  97.39471,
  53.10952,
  96.53465,
  53.65542,
  96.28519,
  53.97191,
  96.77134,
  53.6995,
  97.13009,
  53.30853,
  96.24915,
  53.84383,
  96.13412,
  54.16755,
  96.64586,
  53.82019,
  97.08936,
  53.39629,
  96.4371,
  53.83921,
  95.99113,
  54.13032,
  96.53549,
  53.95083,
  96.90091,
  53.62335,
  96.81501,
  53.55672,
  95.97681,
  54.05401,
  96.26982,
  54.08004,
  75.51859,
  -54.08709,
  75.23147,
  -54.5355,
  75.3961,
  -53.29797,
  75.55688,
  -53.68099,
  75.3566,
  -54.16922,
  75.26958,
  -54.45105,
  75.4162,
  -53.70248,
  75.38531,
  -54.14769,
  75.52645,
  -53.97329,
  75.34688,
  -54.61319,
  75.23702,
  -54.47147,
  75.20194,
  -55.06744,
  75.36372,
  -54.13785,
  75.45895,
  -54.3775,
  75.20199,
  -55.05239,
  75.33098,
  -53.94096,
  75.4597,
  -53.67615,
  75.36191,
  -54.39209,
  75.16953,
  -54.46145,
  75.36732,
  -54.21752,
  75.38213,
  -53.81436,
  75.37733,
  -54.05695,
  75.51015,
  -53.27807,
  75.45236,
  -53.79033,
  75.41233,
  -54.46706,
  75.37808,
  -54.19176,
  75.39451,
  -54.33945,
  75.39181,
  -54.1788,
  75.21043,
  -55.0731,
  75.40028,
  -53.98528,
  75.33826,
  -54.54152,
  75.25341,
  -55.15313,
  75.26748,
  -54.50189,
  75.55816,
  -53.80283,
  75.42896,
  -54.3552,
  75.16218,
  -54.35055,
  75.51836,
  -53.24767,
  75.4175,
  -53.84812,
  75.55477,
  -54.16561,
  75.42219,
  -53.66631,
  75.54333,
  -53.46295,
  75.58223,
  -53.52993,
  75.49554,
  -53.94402,
  75.32068,
  -54.61244,
  75.22739,
  -54.98266,
  75.21947,
  -54.63861,
  75.41308,
  -54.04442,
  75.45478,
  -54.39002,
  75.27288,
  -55.04627,
  75.12544,
  -55.18523,
  75.32343,
  -53.80637,
  75.39137,
  -54.30791,
  75.38635,
  -54.82091,
  75.21485,
  -54.68422,
  75.56799,
  -53.4447,
  75.61134,
  -53.93412,
  75.2687,
  -54.47602,
  75.34281,
  -53.5691,
  75.4961,
  -53.82009,
  75.39876,
  -53.8718,
  75.44255,
  -54.09045,
  75.41682,
  -54.20765,
  75.25925,
  -54.52288,
  75.31283,
  -53.82047,
  75.53893,
  -54.13307,
  75.31055,
  -54.48671,
  75.26873,
  -54.86162,
  75.35027,
  -54.76934,
  75.38833,
  -54.34781,
  75.36046,
  -54.65005,
  75.21769,
  -55.18739,
  75.20079,
  -54.65434,
  75.52124,
  -53.78849,
  75.31606,
  -54.48901,
  75.19054,
  -55.03466,
  75.32172,
  -53.92942,
  75.42559,
  -53.61789,
  75.33719,
  -54.26687,
  75.31184,
  -54.72097,
  75.32565,
  -53.86648,
  75.34958,
  -53.54819,
  75.46464,
  -54.10466,
  75.37309,
  -54.57225,
  75.31036,
  -54.39969,
  75.398,
  -53.56993,
  75.52962,
  -53.83891,
  75.44175,
  -53.93009,
  75.22988,
  -54.75896,
  75.17886,
  -54.80185,
  75.43018,
  -53.98878,
  75.42763,
  -54.18171,
  75.45654,
  -54.48278,
  75.26601,
  -55.15636,
  75.34913,
  -54.569,
  75.46776,
  -54.19893,
  75.3456,
  -54.75824,
  75.26219,
  -55.2667,
  75.23088,
  -54.58926,
  75.41037,
  -53.88054,
  75.50363,
  -54.37549,
  75.33134,
  -54.99093,
  75.26569,
  -54.39549,
  75.55569,
  -53.57841,
  75.5463,
  -54.2833,
  75.25081,
  -54.89548,
  75.41616,
  -53.79699,
  75.45458,
  -53.53382,
  75.39362,
  -54.10411,
  75.33014,
  -54.58737,
  75.35191,
  -54.41789,
  75.41148,
  -53.51297,
  75.43633,
  -53.90536,
  75.46191,
  -54.22391,
  75.49309,
  -54.52798,
  75.20796,
  -54.40123,
  75.43697,
  -53.60555,
  75.52506,
  -54.13408,
  75.33442,
  -54.64255,
  75.13214,
  -55.10266,
  75.18999,
  -54.40135,
  75.43524,
  -53.96434,
  75.26932,
  -54.18369,
  75.21095,
  -55.11829,
  75.13557,
  -55.37659,
  75.2363,
  -54.49734,
  75.41742,
  -54.48114,
  75.28939,
  -54.89066,
  75.1829,
  -55.10565,
  75.24188,
  -53.90519,
  75.52155,
  -54.08765,
  75.38099,
  -54.68324,
  75.08833,
  -55.16176,
  75.1459,
  -53.908,
  75.53945,
  -53.85357,
  75.35417,
  -54.55063,
  75.12238,
  -55.02716,
  75.30126,
  -54.11128,
  75.50228,
  -53.62773,
  75.39213,
  -54.24347,
  75.28555,
  -54.78887,
  75.28171,
  -53.92458,
  75.43966,
  -53.57539,
  75.47146,
  -53.9573,
  75.3376,
  -54.44309,
  75.46003,
  -53.50657,
  75.53117,
  -53.32923,
  75.49357,
  -53.80397,
  75.43829,
  -54.30436,
  75.31378,
  -54.77874,
  75.24023,
  -54.13256,
  75.52933,
  -53.80793,
  75.47945,
  -54.37497,
  75.39733,
  -54.57701,
  75.32053,
  -54.77999,
  75.34427,
  -54.1715,
  75.57262,
  -53.81448,
  75.43783,
  -54.56,
  75.28275,
  -55.18037,
  75.23969,
  -55.55927,
  75.50911,
  -54.37379,
  75.41422,
  -54.41987,
  75.34859,
  -54.86227,
  75.16001,
  -55.3903,
  75.21913,
  -54.26826,
  75.53616,
  -54.10493,
  75.39699,
  -54.67525,
  75.1858,
  -55.14968,
  75.42086,
  -54.06858,
  75.59429,
  -53.76233,
  75.31252,
  -54.48466,
  75.28884,
  -55.01132,
  75.30601,
  -53.95227,
  75.41367,
  -53.64331,
  75.37709,
  -54.16016,
  75.40265,
  -54.49108,
  75.405,
  -53.29064,
  75.43598,
  -53.27973,
  75.55351,
  -53.97705,
  75.35275,
  -54.53227,
  75.26194,
  -54.41441,
  75.51382,
  -53.25823,
  75.53917,
  -53.67912,
  75.32951,
  -54.31174,
  75.39924,
  -54.6587,
  75.35934,
  -53.83406,
  75.42509,
  -53.57505,
  75.42735,
  -54.31968,
  75.50877,
  -54.77357,
  75.3229,
  -54.737,
  75.36761,
  -53.98958,
  75.47401,
  -53.83375,
  75.48244,
  -54.4837,
  75.22174,
  -54.77822,
  75.22047,
  -54.5752,
  75.49251,
  -53.80748,
  75.44043,
  -54.33756,
  75.3713,
  -54.68293,
  75.08734,
  -54.84767,
  75.24926,
  -54.74097,
  75.44522,
  -54.16355,
  75.34815,
  -54.69554,
  75.20778,
  -55.18597,
  75.26942,
  -55.25907,
  75.41686,
  -53.98673,
  75.40319,
  -54.46646,
  75.33168,
  -54.97514,
  75.22417,
  -55.08517,
  75.30054,
  -53.92952,
  75.52354,
  -54.14849,
  75.46046,
  -54.74057,
  75.25597,
  -55.12278,
  75.2781,
  -53.70147,
  75.4632,
  -53.84176,
  75.36569,
  -54.47032,
  75.2555,
  -54.80178,
  75.48221,
  -53.31939,
  75.5262,
  -53.7253,
  75.52844,
  -54.26201,
  75.19355,
  -54.77756,
  75.31026,
  -53.63806,
  75.36691,
  -53.46946,
  75.58596,
  -54.0078,
  75.29647,
  -54.51898,
  75.21104,
  -54.4077,
  75.48537,
  -53.46729,
  75.5023,
  -53.93951,
  75.20886,
  -54.46327,
  75.17556,
  -54.51845,
  75.37657,
  -54.26071,
  75.47525,
  -53.72545,
  75.39117,
  -54.21247,
  75.39406,
  -54.56694,
  75.30214,
  -54.39057,
  75.18605,
  -53.80988,
  75.24158,
  -54.45673,
  75.28667,
  -54.56109,
  75.21368,
  -54.58276,
  75.33286,
  -54.18266,
  75.40226,
  -54.24049,
  75.3411,
  -54.38681,
  75.25465,
  -54.84959,
  75.22734,
  -54.39397,
  75.41729,
  -54.11338,
  75.43217,
  -54.14319,
  75.33526,
  -54.74945,
  75.18126,
  -55.28876,
  75.25134,
  -54.3506,
  75.33007,
  -54.06221,
  75.38367,
  -54.58786,
  75.22655,
  -55.14116,
  75.26866,
  -55.26443,
  75.30442,
  -54.03084,
  75.50806,
  -54.10094,
  75.31098,
  -54.76185,
  75.16203,
  -55.2462,
  75.34579,
  -53.96214,
  75.44284,
  -54.07473,
  75.23129,
  -54.55927,
  75.16217,
  -54.91403,
  75.24778,
  -53.61563,
  75.38491,
  -53.64509,
  75.37368,
  -54.47743,
  75.45118,
  -54.93583,
  75.39223,
  -54.15773,
  75.44263,
  -53.53554,
  75.28578,
  -54.05236,
  75.4323,
  -54.61211,
  75.42654,
  -53.9291,
  75.43514,
  -53.67169,
  75.35548,
  -54.11614,
  75.31292,
  -54.33876,
  75.3387,
  -54.20326,
  75.29365,
  -53.43858,
  75.39999,
  -53.57924,
  75.36909,
  -54.14893,
  75.17276,
  -54.76834,
  75.34224,
  -53.64019,
  75.50484,
  -53.60596,
  75.24625,
  -54.56942,
  75.22095,
  -54.61148,
  75.29385,
  -54.72705,
  75.19127,
  -53.99551,
  75.44002,
  -53.89434,
  75.44141,
  -54.35485,
  75.31389,
  -54.74089,
  75.25904,
  -54.57575,
  75.29982,
  -54.36477,
  75.38258,
  -54.33023,
  75.30313,
  -54.6627,
  75.30887,
  -55.04218,
  75.32429,
  -54.72547,
  75.35476,
  -54.17981,
  75.45914,
  -54.28037,
  75.26644,
  -54.76948,
  75.32586,
  -54.67377,
  75.32284,
  -54.19804,
  75.55959,
  -54.1589,
  75.37524,
  -54.78408,
  75.14333,
  -55.13877,
  75.43851,
  -54.02288,
  75.42819,
  -53.97285,
  75.37698,
  -54.48059,
  75.22236,
  -55.08588,
  75.17551,
  -54.0709,
  75.4743,
  -53.68643,
  75.38226,
  -54.37297,
  75.28922,
  -54.82468,
  75.25927,
  -53.79391,
  75.55649,
  -53.5075,
  75.41096,
  -54.07007,
  75.29647,
  -54.62543,
  75.42217,
  -53.9098,
  75.396,
  -53.40115,
  75.4903,
  -53.859,
  75.4784,
  -54.4495,
  75.27647,
  -54.44284,
  75.33399,
  -53.40657,
  75.42719,
  -53.66221,
  -14.22611,
  -77.68449,
  -14.66727,
  -77.65236,
  -13.57793,
  -77.18984,
  -13.94214,
  -77.56248,
  -14.28421,
  -77.55075,
  -14.55616,
  -77.62982,
  -13.86991,
  -77.3364,
  -14.3271,
  -77.6385,
  -14.1154,
  -77.65112,
  -14.71269,
  -77.76078,
  -14.50649,
  -77.6638,
  -15.17249,
  -77.89623,
  -14.32831,
  -77.50005,
  -14.4868,
  -77.81565,
  -15.17351,
  -77.88645,
  -14.14832,
  -77.3691,
  -13.79397,
  -77.50333,
  -14.49368,
  -77.65751,
  -14.60266,
  -77.56497,
  -14.22078,
  -77.4825,
  -14.13271,
  -77.4537,
  -14.19472,
  -77.50739,
  -13.48724,
  -77.26214,
  -13.9379,
  -77.49413,
  -14.61808,
  -77.79191,
  -14.32246,
  -77.56191,
  -14.49095,
  -77.58853,
  -14.36612,
  -77.58026,
  -15.19823,
  -77.77856,
  -14.2,
  -77.51107,
  -14.62934,
  -77.712,
  -15.2589,
  -77.90833,
  -14.69009,
  -77.63795,
  -13.94278,
  -77.59393,
  -14.48192,
  -77.76381,
  -14.64612,
  -77.52103,
  -13.46911,
  -77.20545,
  -14.03464,
  -77.48817,
  -14.25383,
  -77.70805,
  -13.82867,
  -77.36057,
  -13.73678,
  -77.40066,
  -13.68545,
  -77.42338,
  -14.20706,
  -77.59487,
  -14.71686,
  -77.68497,
  -15.03693,
  -77.81213,
  -14.88661,
  -77.71411,
  -14.27692,
  -77.53953,
  -14.50965,
  -77.7781,
  -15.20689,
  -77.85256,
  -15.36814,
  -77.85546,
  -14.05969,
  -77.3513,
  -14.45578,
  -77.6188,
  -14.98228,
  -77.86124,
  -14.94745,
  -77.72793,
  -13.68428,
  -77.42947,
  -14.15347,
  -77.69764,
  -14.79527,
  -77.68385,
  -13.89116,
  -77.29482,
  -14.10654,
  -77.5601,
  -14.09988,
  -77.52631,
  -14.22511,
  -77.61697,
  -14.33797,
  -77.69594,
  -14.71953,
  -77.63065,
  -14.16238,
  -77.39089,
  -14.30371,
  -77.75222,
  -14.65292,
  -77.67383,
  -14.97735,
  -77.82304,
  -14.85907,
  -77.86018,
  -14.52167,
  -77.61987,
  -14.76522,
  -77.79738,
  -15.35681,
  -77.97124,
  -14.94682,
  -77.64253,
  -13.9871,
  -77.60714,
  -14.62699,
  -77.7142,
  -15.19583,
  -77.9387,
  -14.1533,
  -77.34686,
  -13.88076,
  -77.42064,
  -14.46014,
  -77.60462,
  -14.87263,
  -77.77522,
  -14.03466,
  -77.41019,
  -13.83355,
  -77.31379,
  -14.2051,
  -77.65916,
  -14.67204,
  -77.87844,
  -14.529,
  -77.55229,
  -13.78591,
  -77.29118,
  -13.90053,
  -77.56076,
  -14.06005,
  -77.52517,
  -14.85007,
  -77.77479,
  -14.98165,
  -77.68703,
  -14.15705,
  -77.4623,
  -14.35436,
  -77.60439,
  -14.68948,
  -77.7961,
  -15.33887,
  -77.95439,
  -14.74068,
  -77.68169,
  -14.34758,
  -77.67397,
  -14.88284,
  -77.8671,
  -15.39357,
  -78.03759,
  -14.77388,
  -77.63039,
  -14.06666,
  -77.41568,
  -14.55172,
  -77.74725,
  -15.18549,
  -77.8911,
  -14.72207,
  -77.53986,
  -13.88165,
  -77.46487,
  -14.35905,
  -77.72398,
  -14.98699,
  -77.80529,
  -14.03429,
  -77.37096,
  -13.6721,
  -77.33815,
  -14.23597,
  -77.59033,
  -14.70746,
  -77.81149,
  -14.63099,
  -77.71947,
  -13.76768,
  -77.33231,
  -14.0347,
  -77.5126,
  -14.47381,
  -77.71764,
  -14.72417,
  -77.72462,
  -14.50563,
  -77.55444,
  -13.8311,
  -77.45905,
  -14.2625,
  -77.67675,
  -14.89499,
  -77.74629,
  -15.30678,
  -77.8987,
  -14.57711,
  -77.58272,
  -14.12513,
  -77.57543,
  -14.47426,
  -77.56287,
  -15.27161,
  -77.95246,
  -15.57284,
  -77.92033,
  -14.71881,
  -77.59734,
  -14.54914,
  -77.74187,
  -14.91743,
  -77.84224,
  -15.13446,
  -77.93935,
  -14.18128,
  -77.34209,
  -14.29475,
  -77.65765,
  -14.76143,
  -77.8592,
  -15.39743,
  -77.81184,
  -14.17025,
  -77.28748,
  -13.96128,
  -77.50477,
  -14.63412,
  -77.68224,
  -15.16452,
  -77.76639,
  -14.32976,
  -77.42674,
  -13.90117,
  -77.40836,
  -14.42609,
  -77.55147,
  -14.97586,
  -77.78011,
  -14.16573,
  -77.35449,
  -13.83263,
  -77.34474,
  -14.15437,
  -77.56757,
  -14.67096,
  -77.66588,
  -13.72817,
  -77.2532,
  -13.52717,
  -77.27648,
  -14.05219,
  -77.62422,
  -14.45814,
  -77.7288,
  -14.99055,
  -77.82172,
  -14.38631,
  -77.51278,
  -13.89222,
  -77.52826,
  -14.48354,
  -77.72324,
  -14.6524,
  -77.7233,
  -14.88101,
  -77.78097,
  -14.3807,
  -77.58812,
  -14.02726,
  -77.54978,
  -14.64667,
  -77.83348,
  -15.29493,
  -77.97856,
  -15.64287,
  -77.92805,
  -14.54764,
  -77.61349,
  -14.56869,
  -77.71014,
  -14.97384,
  -77.92414,
  -15.43881,
  -77.96307,
  -14.48502,
  -77.47847,
  -14.21796,
  -77.71436,
  -14.73209,
  -77.79946,
  -15.2102,
  -77.9033,
  -14.23137,
  -77.52467,
  -13.80445,
  -77.62361,
  -14.64684,
  -77.71798,
  -15.16628,
  -77.83173,
  -14.16367,
  -77.36317,
  -13.85869,
  -77.29453,
  -14.36021,
  -77.61031,
  -14.71011,
  -77.79643,
  -13.58733,
  -77.2123,
  -13.65087,
  -77.25578,
  -14.11759,
  -77.61141,
  -14.64799,
  -77.82405,
  -14.622,
  -77.59319,
  -13.50153,
  -77.2692,
  -13.92234,
  -77.46346,
  -14.50523,
  -77.64779,
  -14.79593,
  -77.80107,
  -14.06598,
  -77.4876,
  -13.87332,
  -77.30879,
  -14.51872,
  -77.74992,
  -14.85273,
  -77.82487,
  -14.85309,
  -77.7072,
  -14.29099,
  -77.51287,
  -14.07456,
  -77.54951,
  -14.57912,
  -77.77957,
  -14.96981,
  -77.73344,
  -14.83262,
  -77.56297,
  -14.06875,
  -77.49812,
  -14.50031,
  -77.6908,
  -14.79816,
  -77.83287,
  -15.01328,
  -77.65139,
  -14.93933,
  -77.67889,
  -14.29445,
  -77.62045,
  -14.86765,
  -77.74445,
  -15.31992,
  -77.95836,
  -15.39163,
  -78.01579,
  -14.15027,
  -77.52728,
  -14.59214,
  -77.74561,
  -15.10115,
  -77.94356,
  -15.29973,
  -77.87025,
  -14.16257,
  -77.36768,
  -14.26119,
  -77.71517,
  -14.85956,
  -77.93626,
  -15.26915,
  -77.76627,
  -13.97507,
  -77.28825,
  -14.02236,
  -77.61825,
  -14.66078,
  -77.70556,
  -14.9743,
  -77.74224,
  -13.45524,
  -77.28119,
  -13.93555,
  -77.56461,
  -14.50039,
  -77.65386,
  -14.95632,
  -77.80871,
  -13.93687,
  -77.32011,
  -13.80009,
  -77.21938,
  -14.18596,
  -77.72627,
  -14.68249,
  -77.78151,
  -14.6285,
  -77.60478,
  -13.71599,
  -77.29681,
  -14.06586,
  -77.55463,
  -14.62166,
  -77.66806,
  -14.74049,
  -77.78249,
  -14.4505,
  -77.59968,
  -13.93995,
  -77.41051,
  -14.33845,
  -77.60042,
  -14.80618,
  -77.75087,
  -14.65256,
  -77.62537,
  -14.11147,
  -77.25368,
  -14.48204,
  -77.64352,
  -14.71348,
  -77.6834,
  -14.81606,
  -77.6571,
  -14.46154,
  -77.58753,
  -14.42583,
  -77.55718,
  -14.67533,
  -77.58926,
  -15.00728,
  -77.7762,
  -14.58295,
  -77.68156,
  -14.32835,
  -77.58721,
  -14.28408,
  -77.65067,
  -14.89589,
  -77.79637,
  -15.31974,
  -77.90044,
  -14.47767,
  -77.5695,
  -14.22492,
  -77.48806,
  -14.74257,
  -77.61623,
  -15.30886,
  -78.04389,
  -15.23856,
  -77.95309,
  -14.14418,
  -77.48399,
  -14.26879,
  -77.66641,
  -15.11452,
  -77.74654,
  -15.46572,
  -77.95094,
  -14.18366,
  -77.45116,
  -14.20384,
  -77.67905,
  -14.82109,
  -77.66947,
  -15.12344,
  -77.76174,
  -13.94865,
  -77.20683,
  -13.93399,
  -77.41659,
  -14.55163,
  -77.75021,
  -14.96032,
  -77.96703,
  -14.32241,
  -77.55685,
  -13.81945,
  -77.32147,
  -14.33341,
  -77.57384,
  -14.70792,
  -77.71756,
  -14.35042,
  -77.52592,
  -13.83475,
  -77.29808,
  -14.32437,
  -77.54939,
  -14.55144,
  -77.60152,
  -14.44692,
  -77.53131,
  -13.6795,
  -77.15056,
  -13.8709,
  -77.41315,
  -14.29999,
  -77.67805,
  -14.91482,
  -77.78239,
  -13.85426,
  -77.31986,
  -13.80914,
  -77.38786,
  -14.77996,
  -77.66796,
  -14.80933,
  -77.6172,
  -14.92895,
  -77.78773,
  -14.31943,
  -77.33208,
  -14.05001,
  -77.44673,
  -14.53109,
  -77.75127,
  -14.89514,
  -77.86423,
  -14.77049,
  -77.71277,
  -14.60507,
  -77.62816,
  -14.50844,
  -77.65356,
  -14.8162,
  -77.79929,
  -15.16681,
  -77.96514,
  -14.86382,
  -77.75005,
  -14.30791,
  -77.54717,
  -14.44137,
  -77.74139,
  -14.88562,
  -77.82546,
  -14.82699,
  -77.80572,
  -14.35464,
  -77.42073,
  -14.16449,
  -77.68037,
  -14.85523,
  -77.87627,
  -15.28118,
  -77.91873,
  -14.1748,
  -77.55824,
  -14.13898,
  -77.56207,
  -14.68475,
  -77.75585,
  -15.26102,
  -77.82855,
  -14.34724,
  -77.35941,
  -13.91392,
  -77.42021,
  -14.44816,
  -77.67558,
  -14.95393,
  -77.77574,
  -14.07017,
  -77.24312,
  -13.68025,
  -77.39658,
  -14.23736,
  -77.60903,
  -14.87104,
  -77.78573,
  -14.11498,
  -77.42229,
  -13.64874,
  -77.22375,
  -14.03749,
  -77.54807,
  -14.53753,
  -77.74079,
  -14.62295,
  -77.64018,
  -13.69655,
  -77.15564,
  -13.89584,
  -77.37731,
  -65.4136,
  -17.31545,
  -65.66879,
  -16.86457,
  -64.67429,
  -17.64606,
  -65.14156,
  -17.5406,
  -65.36923,
  -17.17989,
  -65.61687,
  -17.00402,
  -65.02346,
  -17.5443,
  -65.43049,
  -17.22604,
  -65.31678,
  -17.40587,
  -65.79259,
  -16.89435,
  -65.51939,
  -16.99392,
  -65.98582,
  -16.56401,
  -65.34724,
  -17.16081,
  -65.67336,
  -17.17053,
  -66.09493,
  -16.52214,
  -65.15239,
  -17.22781,
  -65.13319,
  -17.62809,
  -65.6367,
  -17.1291,
  -65.59461,
  -16.98622,
  -65.24038,
  -17.12525,
  -65.07199,
  -17.30094,
  -65.36268,
  -17.26891,
  -64.68094,
  -17.76766,
  -65.16306,
  -17.4185,
  -65.70817,
  -17.05151,
  -65.54395,
  -17.2228,
  -65.47012,
  -17.04599,
  -65.41509,
  -17.21678,
  -66.05148,
  -16.53701,
  -65.28555,
  -17.37264,
  -65.72754,
  -17.06043,
  -66.15897,
  -16.55838,
  -65.54787,
  -16.95716,
  -65.16622,
  -17.54364,
  -65.59259,
  -17.11258,
  -65.53957,
  -16.87813,
  -64.5818,
  -17.73322,
  -65.1082,
  -17.45738,
  -65.42698,
  -17.35717,
  -64.91531,
  -17.51686,
  -64.94831,
  -17.64612,
  -64.97105,
  -17.69325,
  -65.29108,
  -17.33554,
  -65.73941,
  -16.9185,
  -66.02723,
  -16.57476,
  -65.69793,
  -16.80672,
  -65.35004,
  -17.24775,
  -65.71232,
  -17.19592,
  -66.14458,
  -16.64243,
  -66.08742,
  -16.45742,
  -65.05412,
  -17.3876,
  -65.50035,
  -17.14974,
  -65.8932,
  -16.8185,
  -65.66531,
  -16.77991,
  -64.91454,
  -17.70176,
  -65.36417,
  -17.4383,
  -65.65968,
  -16.928,
  -64.92522,
  -17.45603,
  -65.16066,
  -17.36914,
  -65.17289,
  -17.37957,
  -65.29445,
  -17.31087,
  -65.42591,
  -17.24259,
  -65.59834,
  -16.90846,
  -65.0518,
  -17.31906,
  -65.56509,
  -17.27248,
  -65.61161,
  -17.02073,
  -65.80602,
  -16.7756,
  -65.84576,
  -16.85386,
  -65.48976,
  -17.15793,
  -65.77794,
  -16.94801,
  -66.22222,
  -16.54594,
  -65.69975,
  -16.7118,
  -65.19217,
  -17.52367,
  -65.71246,
  -16.99064,
  -66.14365,
  -16.56097,
  -65.0961,
  -17.25074,
  -65.07049,
  -17.52748,
  -65.53711,
  -17.12208,
  -65.84769,
  -16.78749,
  -65.13745,
  -17.24428,
  -64.8541,
  -17.46768,
  -65.49252,
  -17.34868,
  -65.80704,
  -17.07225,
  -65.47779,
  -17.06184,
  -64.90906,
  -17.62169,
  -65.36239,
  -17.52216,
  -65.23944,
  -17.36934,
  -65.87533,
  -16.86575,
  -65.79723,
  -16.68737,
  -65.25683,
  -17.29705,
  -65.45023,
  -17.19605,
  -65.73119,
  -17.16815,
  -66.20834,
  -16.48936,
  -65.63289,
  -16.90127,
  -65.43767,
  -17.21124,
  -65.80921,
  -16.85065,
  -66.26577,
  -16.50797,
  -65.65154,
  -16.7652,
  -65.15229,
  -17.35793,
  -65.58071,
  -17.05051,
  -66.06771,
  -16.62245,
  -65.4465,
  -16.88117,
  -64.9891,
  -17.56809,
  -65.56495,
  -17.24459,
  -65.89011,
  -16.73516,
  -65.03742,
  -17.44224,
  -64.84667,
  -17.79194,
  -65.36618,
  -17.33582,
  -65.87181,
  -16.91163,
  -65.6152,
  -17.01048,
  -64.80544,
  -17.53041,
  -65.11933,
  -17.39159,
  -65.54987,
  -17.14266,
  -65.67567,
  -16.93864,
  -65.4463,
  -16.9363,
  -65.06026,
  -17.50682,
  -65.5189,
  -17.29402,
  -65.80636,
  -16.91574,
  -66.06483,
  -16.49912,
  -65.53575,
  -16.92817,
  -65.28113,
  -17.32918,
  -65.53261,
  -17.1174,
  -66.21879,
  -16.63403,
  -66.34425,
  -16.27964,
  -65.66501,
  -16.93845,
  -65.56926,
  -16.97583,
  -65.939,
  -16.7079,
  -66.02677,
  -16.57191,
  -65.04559,
  -17.21778,
  -65.2891,
  -17.36287,
  -65.80398,
  -16.94683,
  -66.14074,
  -16.37448,
  -65.06702,
  -17.1872,
  -65.23199,
  -17.50333,
  -65.60998,
  -16.99762,
  -65.93317,
  -16.53249,
  -65.19358,
  -17.09374,
  -64.98878,
  -17.56582,
  -65.48833,
  -17.18112,
  -65.8596,
  -16.7384,
  -65.14354,
  -17.21918,
  -64.92284,
  -17.56188,
  -65.30698,
  -17.29184,
  -65.71272,
  -16.96788,
  -64.85424,
  -17.57573,
  -64.69997,
  -17.73363,
  -65.25862,
  -17.49399,
  -65.59097,
  -17.1166,
  -65.8697,
  -16.82237,
  -65.3186,
  -17.10605,
  -65.13284,
  -17.50175,
  -65.52362,
  -17.20177,
  -65.71736,
  -17.0102,
  -65.81969,
  -16.768,
  -65.38956,
  -17.11209,
  -65.3202,
  -17.45334,
  -65.73111,
  -17.02074,
  -66.14649,
  -16.61606,
  -66.36336,
  -16.35251,
  -65.61518,
  -17.09956,
  -65.63387,
  -17.04305,
  -65.99941,
  -16.87428,
  -66.25779,
  -16.43367,
  -65.32607,
  -16.94483,
  -65.28927,
  -17.28366,
  -65.8113,
  -16.87819,
  -66.07552,
  -16.55594,
  -65.25752,
  -17.32905,
  -65.21776,
  -17.55762,
  -65.68289,
  -17.02563,
  -66.0263,
  -16.67901,
  -65.24593,
  -17.24352,
  -64.99786,
  -17.53933,
  -65.55932,
  -17.20984,
  -65.70011,
  -17.02349,
  -64.72225,
  -17.67297,
  -64.65107,
  -17.69513,
  -65.34717,
  -17.4549,
  -65.70824,
  -17.01204,
  -65.48903,
  -17.00043,
  -64.70119,
  -17.77437,
  -65.11494,
  -17.56878,
  -65.57893,
  -17.06824,
  -65.84303,
  -16.93047,
  -65.15114,
  -17.43583,
  -64.90158,
  -17.55132,
  -65.60751,
  -17.19142,
  -65.93345,
  -16.90702,
  -65.7959,
  -16.84223,
  -65.30917,
  -17.23953,
  -65.19015,
  -17.39762,
  -65.68808,
  -17.07271,
  -65.89011,
  -16.7203,
  -65.73384,
  -16.78081,
  -65.18789,
  -17.4627,
  -65.48322,
  -17.17061,
  -65.89466,
  -16.91747,
  -65.82989,
  -16.70115,
  -65.79685,
  -16.6877,
  -65.43296,
  -17.19184,
  -65.79544,
  -16.84646,
  -66.20834,
  -16.44394,
  -66.25231,
  -16.47211,
  -65.31441,
  -17.30787,
  -65.64532,
  -17.07093,
  -66.04717,
  -16.75897,
  -66.11391,
  -16.5124,
  -65.09577,
  -17.27048,
  -65.42595,
  -17.33057,
  -65.92611,
  -16.88039,
  -66.1107,
  -16.53036,
  -64.94862,
  -17.42986,
  -65.32838,
  -17.54066,
  -65.69572,
  -17.01096,
  -65.92395,
  -16.61395,
  -64.67792,
  -17.71678,
  -65.12124,
  -17.52883,
  -65.52708,
  -17.25541,
  -65.86211,
  -16.82232,
  -64.96172,
  -17.38801,
  -64.81756,
  -17.59214,
  -65.3383,
  -17.36878,
  -65.70287,
  -17.07122,
  -65.52787,
  -16.93734,
  -64.84846,
  -17.66766,
  -65.2864,
  -17.42506,
  -65.63422,
  -17.03601,
  -65.71009,
  -16.79371,
  -65.4334,
  -17.09656,
  -65.0999,
  -17.38993,
  -65.55564,
  -17.21666,
  -65.81474,
  -16.94444,
  -65.5048,
  -17.01373,
  -65.00552,
  -17.33883,
  -65.6601,
  -16.93491,
  -65.66124,
  -16.7982,
  -65.65498,
  -16.75309,
  -65.43763,
  -17.0482,
  -65.52513,
  -17.10456,
  -65.60825,
  -16.98089,
  -65.88806,
  -16.70184,
  -65.47815,
  -16.92927,
  -65.40737,
  -17.12625,
  -65.42101,
  -17.22795,
  -65.81525,
  -16.82844,
  -66.15499,
  -16.46707,
  -65.66698,
  -17.02043,
  -65.22378,
  -17.2444,
  -65.71648,
  -16.90278,
  -66.21609,
  -16.59329,
  -66.2047,
  -16.51548,
  -65.17854,
  -17.28729,
  -65.50632,
  -17.3997,
  -65.96799,
  -16.90122,
  -66.2174,
  -16.42444,
  -65.1788,
  -17.24247,
  -65.43721,
  -17.34045,
  -65.69265,
  -16.82738,
  -65.96646,
  -16.59011,
  -64.84525,
  -17.28774,
  -65.06837,
  -17.49044,
  -65.63849,
  -17.08027,
  -66.04486,
  -16.82393,
  -65.3046,
  -17.20261,
  -64.91376,
  -17.57021,
  -65.43085,
  -17.27434,
  -65.74316,
  -16.83323,
  -65.22941,
  -17.25269,
  -64.91863,
  -17.53299,
  -65.27059,
  -17.20961,
  -65.53589,
  -17.02228,
  -65.45172,
  -17.14399,
  -64.70564,
  -17.53323,
  -64.93234,
  -17.52777,
  -65.40356,
  -17.27291,
  -65.7463,
  -16.81972,
  -64.94446,
  -17.54501,
  -64.9896,
  -17.57903,
  -65.65927,
  -16.86263,
  -65.66424,
  -16.79192,
  -65.85395,
  -16.86788,
  -65.11132,
  -17.14472,
  -65.13326,
  -17.43316,
  -65.6098,
  -17.18105,
  -65.99287,
  -16.81831,
  -65.69089,
  -16.87596,
  -65.55578,
  -17.01327,
  -65.51942,
  -17.11365,
  -65.77191,
  -16.84866,
  -66.03346,
  -16.62074,
  -65.81143,
  -16.80344,
  -65.39483,
  -17.2298,
  -65.56667,
  -17.11049,
  -65.87546,
  -16.78226,
  -65.81636,
  -16.86609,
  -65.26316,
  -17.15839,
  -65.43443,
  -17.31758,
  -65.85508,
  -16.88068,
  -66.06793,
  -16.57218,
  -65.21304,
  -17.31335,
  -65.21503,
  -17.34257,
  -65.70286,
  -17.01162,
  -66.12071,
  -16.57997,
  -65.1683,
  -17.06827,
  -65.10743,
  -17.47272,
  -65.5929,
  -17.11454,
  -65.86874,
  -16.78018,
  -64.96012,
  -17.31385,
  -64.92161,
  -17.65481,
  -65.3351,
  -17.1768,
  -65.81267,
  -16.82844,
  -65.19736,
  -17.30173,
  -64.74113,
  -17.70844,
  -65.2647,
  -17.44154,
  -65.65023,
  -17.07519,
  -65.54909,
  -17.01077,
  -64.68964,
  -17.55024,
  -65.0283,
  -17.5191 ;

 srcpos =
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626244, 5611928, 10.64177, 115.9334, 42.24449, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626300, 5611985, 10.69029, 115.7091, 42.52022, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626355, 5612044, 10.57828, 115.6839, 43.12244, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626411, 5612101, 10.58254, 115.5409, 43.16796, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626468, 5612157, 10.69505, 115.5339, 42.6991, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626525, 5612213, 10.72602, 114.7859, 42.44717, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626581, 5612270, 10.7667, 114.367, 42.24209, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626638, 5612327, 10.7502, 114.5699, 42.0361, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626694, 5612384, 10.66169, 114.6542, 41.61217, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626750, 5612441, 10.56953, 114.9736, 41.33253, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626806, 5612498, 10.57526, 114.9706, 41.35981, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626862, 5612555, 10.67585, 115.7628, 41.27157, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626918, 5612612, 10.7069, 115.5178, 41.3956, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1626973, 5612671, 10.61673, 114.0913, 41.52151, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627027, 5612729, 10.60478, 113.7961, 41.80894, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627082, 5612788, 10.70146, 113.8579, 42.04467, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627137, 5612846, 10.70803, 114.4182, 42.32093, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627192, 5612904, 10.68775, 114.9389, 42.18502, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627246, 5612963, 10.61209, 115.0781, 42.3364, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627300, 5613021, 10.63574, 115.1485, 43.06088, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627355, 5613079, 10.68422, 115.3273, 43.47659, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627410, 5613138, 10.65488, 115.9267, 43.97235, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627465, 5613196, 10.70915, 116.3099, 44.42759, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627520, 5613254, 10.66912, 115.9168, 44.83314, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627575, 5613312, 10.52593, 114.663, 45.54781, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627631, 5613370, 10.50475, 114.8339, 45.81888, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627686, 5613428, 10.5512, 115.8664, 46.08248, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627741, 5613486, 10.61932, 115.8028, 46.62973, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627796, 5613543, 10.69697, 114.6955, 46.78429, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627852, 5613601, 10.6763, 114.6647, 46.95648, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627908, 5613658, 10.5835, 115.1938, 47.06494, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1627964, 5613715, 10.55088, 115.2845, 46.78111, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628020, 5613772, 10.53751, 115.068, 46.70215, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628077, 5613829, 10.60662, 114.7911, 46.31573, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628132, 5613886, 10.60719, 114.8472, 46.22446, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628188, 5613944, 10.54412, 115.199, 46.64112, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628244, 5614000, 10.60878, 114.9755, 47.0546, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628301, 5614057, 10.73807, 115.119, 47.01254, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628359, 5614113, 10.77943, 115.1087, 45.9893, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628416, 5614168, 10.79471, 114.553, 44.62094, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628473, 5614224, 10.85771, 114.4094, 43.83631, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628530, 5614280, 10.87343, 114.8026, 43.27702, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628587, 5614337, 10.89364, 114.4393, 43.15963, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628643, 5614393, 10.89581, 114.0319, 42.72105, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628701, 5614449, 10.87177, 114.1886, 42.35485, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628758, 5614505, 10.93644, 114.2369, 41.77559, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628815, 5614561, 10.90757, 114.468, 41.20041, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628872, 5614617, 10.83352, 114.0639, 40.55069, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628929, 5614674, 10.87408, 114.1099, 39.39336, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1628985, 5614731, 10.8016, 114.5219, 38.5445, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629041, 5614788, 10.76621, 114.5927, 38.73448, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629096, 5614846, 10.79208, 115.2964, 39.1526, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629150, 5614905, 10.73356, 114.6092, 40.15412, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629204, 5614964, 10.68174, 113.219, 40.84945, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629259, 5615023, 10.68063, 113.9009, 41.58089, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629313, 5615082, 10.66602, 114.0638, 42.46506, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629367, 5615140, 10.67172, 113.8734, 43.05365, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629423, 5615198, 10.75093, 114.0892, 43.32463, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629478, 5615256, 10.75049, 114.3524, 43.7948, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629532, 5615314, 10.72055, 114.55, 44.39148, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629587, 5615374, 10.65843, 114.2063, 45.28197, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629641, 5615432, 10.60368, 114.523, 45.71692, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629696, 5615490, 10.63774, 114.4335, 45.77457, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629751, 5615547, 10.58505, 114.0667, 45.58339, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629808, 5615605, 10.58337, 114.4864, 45.66576, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629863, 5615662, 10.57804, 114.8268, 45.73968, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629919, 5615720, 10.54241, 114.4982, 45.82907, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1629975, 5615776, 10.58723, 114.538, 45.71378, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630032, 5615834, 10.61697, 114.3499, 45.53118, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630088, 5615890, 10.64055, 115.1958, 45.47557, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630144, 5615947, 10.65746, 115.3427, 45.35678, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630199, 5616004, 10.59308, 114.7033, 45.19156, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630255, 5616062, 10.62452, 114.4016, 45.51311, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630310, 5616120, 10.66179, 113.8295, 45.64887, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630365, 5616178, 10.66698, 113.7997, 45.48392, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630423, 5616234, 10.66916, 113.8477, 44.78429, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630479, 5616291, 10.6315, 114.4047, 44.24866, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630535, 5616349, 10.66718, 114.509, 44.5905, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630590, 5616406, 10.71402, 114.8471, 45.12468, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630645, 5616464, 10.67367, 114.9045, 45.73659, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630701, 5616521, 10.67033, 114.3212, 45.61581, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630758, 5616578, 10.69564, 113.8055, 44.98746, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630814, 5616635, 10.59346, 114.0768, 44.48682, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630870, 5616693, 10.5479, 114.5529, 44.64349, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630924, 5616750, 10.59712, 115.2108, 44.97446, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1630980, 5616808, 10.60357, 114.7807, 45.16546, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631036, 5616865, 10.5912, 113.9265, 45.22147, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631092, 5616922, 10.63393, 114.0336, 45.08529, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631147, 5616979, 10.61306, 113.648, 45.19523, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631204, 5617038, 10.57333, 113.232, 45.48895, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631259, 5617094, 10.54658, 113.9708, 45.73949, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631316, 5617151, 10.63028, 113.9801, 45.35691, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631372, 5617207, 10.67747, 113.9166, 44.99868, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631429, 5617264, 10.56713, 113.8144, 44.53553, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631485, 5617321, 10.52927, 113.1879, 44.57142, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631541, 5617378, 10.51684, 113.1349, 44.83042, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631597, 5617435, 10.54239, 113.611, 44.85392, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631654, 5617492, 10.59571, 113.7824, 44.51821, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631710, 5617549, 10.60226, 113.6982, 44.27954, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631766, 5617606, 10.61712, 113.8937, 44.3171, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631822, 5617663, 10.69342, 114.076, 43.89642, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631879, 5617720, 10.74287, 113.8797, 43.38466, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631934, 5617778, 10.6673, 113.2008, 43.58861, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1631988, 5617837, 10.58671, 113.2232, 43.90026, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632043, 5617895, 10.59342, 114.2709, 43.90511, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632098, 5617952, 10.58593, 114.5421, 44.06057, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632154, 5618010, 10.53515, 114.1597, 44.04439, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632209, 5618068, 10.57169, 115.0269, 44.42869, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632264, 5618126, 10.60707, 114.7287, 45.14364, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632320, 5618184, 10.49756, 113.6213, 44.95931, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632375, 5618241, 10.46367, 113.5825, 44.97728, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632431, 5618298, 10.60761, 114.3455, 44.95267, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632486, 5618356, 10.62824, 114.7215, 45.27442, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632541, 5618414, 10.60018, 113.8979, 45.53953, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632597, 5618471, 10.66227, 114.0186, 45.82295, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632652, 5618530, 10.65239, 113.8102, 45.97533, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632707, 5618588, 10.65941, 112.9406, 46.63124, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632762, 5618646, 10.64264, 112.69, 47.17958, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632818, 5618703, 10.58387, 113.274, 46.96028, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632873, 5618761, 10.50012, 113.7816, 46.97671, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632929, 5618819, 10.54359, 113.9824, 47.42012, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1632985, 5618876, 10.66836, 114.9286, 47.30351, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633041, 5618932, 10.67659, 114.5217, 47.15397, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633097, 5618989, 10.64312, 112.9023, 46.81959, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633153, 5619046, 10.58815, 113.1633, 46.55078, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633208, 5619105, 10.49634, 114.1431, 46.79524, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633263, 5619163, 10.4858, 114.2861, 47.62718, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633319, 5619220, 10.56072, 114.5459, 47.96753, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633375, 5619278, 10.50536, 114.8216, 48.10231, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633432, 5619334, 10.5387, 113.8908, 47.89457, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633488, 5619390, 10.61163, 114.1364, 46.78909, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633545, 5619447, 10.5994, 114.4818, 46.41337, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633602, 5619504, 10.61696, 114.1521, 46.54292, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633659, 5619559, 10.65582, 114.3902, 46.08749, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633716, 5619616, 10.64665, 113.7801, 45.36877, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633771, 5619673, 10.55566, 112.8623, 44.7845, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633827, 5619731, 10.57882, 112.5644, 45.00196, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633881, 5619789, 10.64452, 112.7501, 45.43541, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633936, 5619848, 10.63358, 112.8048, 46.35847, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1633991, 5619906, 10.55449, 113.2015, 46.82647, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634047, 5619963, 10.53594, 113.7737, 46.53909, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634103, 5620020, 10.55617, 114.3561, 45.87344, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634159, 5620077, 10.59734, 114.7686, 45.80083, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634215, 5620134, 10.56585, 113.9693, 46.42392, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634272, 5620191, 10.58212, 113.4502, 46.5695, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634329, 5620247, 10.62456, 114.4857, 46.24678, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634386, 5620303, 10.62748, 113.6958, 45.51069, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634443, 5620359, 10.65945, 112.8625, 44.51742, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634499, 5620416, 10.67812, 113.1522, 44.39728, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634554, 5620473, 10.66417, 112.8868, 44.98951, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634610, 5620531, 10.628, 112.5506, 44.81084, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634666, 5620588, 10.57455, 113.0152, 44.61887, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634723, 5620646, 10.58369, 113.2092, 44.46714, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634778, 5620703, 10.60047, 112.8119, 44.66912, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634834, 5620760, 10.57833, 113.3178, 44.68589, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634890, 5620816, 10.5826, 113.5302, 44.37594, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1634947, 5620873, 10.56625, 113.0944, 44.0379, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635003, 5620931, 10.62871, 113.1319, 44.08879, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635058, 5620988, 10.65582, 113.359, 44.22656, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635114, 5621045, 10.66588, 112.8472, 44.38095, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635170, 5621102, 10.74117, 112.3519, 44.46178, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635227, 5621159, 10.77052, 112.246, 44.42457, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635283, 5621215, 10.78149, 112.3635, 43.68746, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635339, 5621273, 10.72251, 112.5596, 43.16714, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635394, 5621331, 10.70168, 112.0166, 43.36623, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635449, 5621389, 10.69024, 112.1076, 43.58594, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635503, 5621448, 10.63969, 112.654, 44.81706, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635558, 5621506, 10.68893, 112.5633, 45.65428, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635614, 5621564, 10.68169, 112.1409, 45.93149, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635670, 5621621, 10.64495, 112.3756, 45.40262, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635727, 5621677, 10.63462, 112.3234, 44.80496, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635783, 5621734, 10.62291, 112.0324, 44.1823, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635839, 5621791, 10.6031, 112.3242, 44.00341, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635894, 5621849, 10.59946, 112.627, 44.01666, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1635948, 5621908, 10.6158, 112.2498, 44.77808, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636002, 5621968, 10.66023, 112.4763, 45.63347, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636057, 5622026, 10.69636, 112.6605, 46.26753, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636112, 5622084, 10.66698, 112.6742, 46.70475, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636167, 5622142, 10.55521, 112.6538, 47.16979, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636221, 5622201, 10.50966, 112.2578, 47.73708, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636278, 5622257, 10.57779, 112.2653, 47.8804, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636335, 5622314, 10.5743, 112.2989, 47.72609, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636392, 5622369, 10.56654, 112.3444, 47.28837, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636450, 5622425, 10.6565, 112.6483, 46.21044, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636506, 5622481, 10.70819, 112.7598, 45.45285, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636561, 5622540, 10.60535, 112.1744, 45.32886, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636615, 5622599, 10.59866, 112.4119, 46.24784, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636668, 5622659, 10.61251, 112.6379, 47.43874, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636721, 5622719, 10.68231, 112.9953, 48.93853, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636774, 5622779, 10.69534, 113.3415, 50.24207, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636827, 5622838, 10.6758, 112.7669, 51.05426, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636883, 5622897, 10.71559, 112.9833, 52.07264, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636938, 5622953, 10.64425, 112.8687, 53.22054, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1636995, 5623010, 10.59015, 112.2872, 53.51109, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637053, 5623065, 10.59369, 112.3234, 52.01783, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637111, 5623120, 10.5905, 112.2407, 49.81876, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637169, 5623176, 10.63657, 112.0431, 48.955, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637225, 5623234, 10.65499, 111.9817, 49.11259, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637279, 5623291, 10.62328, 111.7288, 49.43167, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637336, 5623349, 10.57653, 111.6174, 49.22352, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637392, 5623406, 10.59189, 111.5724, 49.09755, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637447, 5623463, 10.56628, 112.4791, 49.37954, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637502, 5623521, 10.5939, 112.2871, 50.04329, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637561, 5623577, 10.58889, 111.7673, 49.51888, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637617, 5623632, 10.43886, 112.4784, 48.63625, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637675, 5623689, 10.49837, 112.5563, 47.68764, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637732, 5623744, 10.55455, 112.4776, 47.20655, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637787, 5623802, 10.3998, 112.0221, 47.39978, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637841, 5623862, 10.38013, 112.5306, 47.46167, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637895, 5623921, 10.4877, 114.2736, 48.07, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1637948, 5623981, 10.49979, 113.4013, 48.74976, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638001, 5624041, 10.50188, 112.5793, 49.7696, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638054, 5624101, 10.59389, 112.9185, 51.3428, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638107, 5624161, 10.61827, 112.4167, 52.83067, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638161, 5624220, 10.65018, 112.6576, 53.86221, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638217, 5624276, 10.57906, 112.3175, 54.86465, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638276, 5624332, 10.49829, 111.7477, 54.8857, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638336, 5624385, 10.56651, 111.8639, 53.20253, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638394, 5624438, 10.59236, 112.3906, 51.57647, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638454, 5624494, 10.62402, 112.3517, 50.99525, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638510, 5624550, 10.58241, 111.8502, 50.6974, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638565, 5624607, 10.64781, 111.8834, 50.48643, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638620, 5624667, 10.71718, 112.549, 51.04068, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638673, 5624727, 10.59947, 112.4561, 52.52609, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638726, 5624786, 10.46667, 111.9061, 54.38118, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638781, 5624844, 10.46541, 112.1607, 54.83128, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638838, 5624900, 10.55082, 112.18, 53.46213, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638894, 5624958, 10.56521, 113.0048, 52.86134, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1638949, 5625016, 10.57316, 112.8207, 53.22892, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639002, 5625076, 10.61259, 112.5167, 54.22021, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639056, 5625135, 10.60519, 112.4437, 55.39445, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639109, 5625194, 10.59131, 111.874, 57.14101, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639165, 5625252, 10.61161, 112.398, 58.20173, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639223, 5625307, 10.62544, 112.2218, 57.69516, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639283, 5625361, 10.60423, 111.2934, 56.83068, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639341, 5625416, 10.53831, 111.8353, 56.17993, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639399, 5625471, 10.55428, 112.4706, 55.94182, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639456, 5625528, 10.65649, 112.3673, 55.87586, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639511, 5625585, 10.63056, 112.8335, 56.01137, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639567, 5625642, 10.59504, 112.5952, 56.4568, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639623, 5625699, 10.5838, 111.8102, 56.72184, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639682, 5625754, 10.58205, 112.1879, 55.98352, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639741, 5625808, 10.52153, 113.8472, 54.64717, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639800, 5625863, 10.55159, 115.1406, 53.57976, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639858, 5625918, 10.61995, 113.0945, 52.23376, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639915, 5625974, 10.57559, 111.1704, 50.73646, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1639970, 5626032, 10.56923, 112.1227, 49.69291, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640022, 5626093, 10.60724, 112.9247, 50.23892, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640073, 5626154, 10.58124, 112.3845, 51.42928, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640124, 5626217, 10.4255, 111.6202, 53.96526, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640176, 5626278, 10.41352, 112.5369, 57.27967, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640231, 5626336, 10.50356, 113.4155, 59.10028, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640287, 5626392, 10.48364, 111.5413, 59.54842, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640346, 5626447, 10.50142, 110.9856, 58.82182, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640405, 5626502, 10.60479, 112.4441, 57.10591, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640461, 5626558, 10.70823, 111.846, 55.93587, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640516, 5626617, 10.64696, 110.4841, 56.04365, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640568, 5626678, 10.54781, 110.9524, 56.49495, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640619, 5626739, 10.56166, 111.1964, 57.81924, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640671, 5626800, 10.59791, 111.5677, 60.0034, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640724, 5626861, 10.58034, 112.6301, 61.34895, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640779, 5626918, 10.61608, 111.9428, 62.44268, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640837, 5626974, 10.5722, 110.6376, 62.07367, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640895, 5627029, 10.56988, 111.1642, 60.69328, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1640952, 5627085, 10.54613, 111.2815, 59.36523, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641009, 5627142, 10.609, 111.6581, 59.18212, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641065, 5627198, 10.67377, 111.8037, 59.84315, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641124, 5627252, 10.55342, 112.3693, 60.67446, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641184, 5627305, 10.48969, 112.1235, 61.07744, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641244, 5627359, 10.521, 111.734, 59.64781, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641303, 5627413, 10.64535, 111.2537, 58.27758, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641359, 5627471, 10.61498, 111.2379, 57.08702, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641412, 5627531, 10.62014, 111.6176, 57.52055, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641466, 5627590, 10.72191, 111.0494, 58.44759, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641520, 5627648, 10.69521, 110.5704, 58.45173, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641577, 5627706, 10.64158, 110.882, 58.42231, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641633, 5627762, 10.57098, 111.0996, 58.66461, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641689, 5627819, 10.59568, 110.8542, 58.32594, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641746, 5627876, 10.62503, 110.9888, 57.83797, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641802, 5627933, 10.54909, 111.3854, 58.10649, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641856, 5627991, 10.53827, 111.6406, 58.58986, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641910, 5628050, 10.52578, 112.4692, 58.87067, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1641965, 5628108, 10.56488, 111.8672, 59.54456, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642022, 5628165, 10.59645, 111.1395, 59.68547, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642079, 5628221, 10.62024, 111.6384, 59.32601, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642137, 5628277, 10.56444, 111.4106, 58.41234, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642195, 5628332, 10.49289, 111.6014, 57.46619, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642253, 5628386, 10.50839, 111.3999, 56.1099, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642310, 5628443, 10.45778, 111.4198, 55.57929, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642365, 5628502, 10.42385, 111.8895, 55.11609, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642418, 5628560, 10.42661, 111.4689, 55.71194, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642472, 5628620, 10.43063, 112.2699, 56.75195, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642527, 5628678, 10.46004, 112.297, 57.24702, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642581, 5628736, 10.54463, 111.2378, 57.47275, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642637, 5628795, 10.53531, 110.9932, 57.76483, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642691, 5628853, 10.40921, 111.0354, 58.61037, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642745, 5628912, 10.39055, 112.4651, 59.82129, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642800, 5628971, 10.371, 112.846, 60.57578, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642856, 5629028, 10.43739, 111.673, 60.42466, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642912, 5629084, 10.47481, 111.8597, 59.91111, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1642968, 5629143, 10.42326, 112.3335, 60.25059, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643022, 5629200, 10.44881, 111.0464, 60.97358, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643079, 5629258, 10.54578, 110.9686, 60.61148, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643135, 5629314, 10.54475, 111.9271, 60.05669, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643192, 5629371, 10.55317, 111.6027, 59.55702, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643248, 5629427, 10.54568, 111.8135, 59.0892, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643305, 5629485, 10.48361, 112.5757, 58.79021, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643362, 5629540, 10.46239, 112.7177, 58.61145, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643419, 5629597, 10.44038, 112.4846, 58.27707, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643476, 5629653, 10.39519, 112.3778, 57.36971, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643533, 5629708, 10.39496, 112.4726, 56.45069, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643590, 5629765, 10.46615, 111.5495, 55.98907, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643647, 5629821, 10.44483, 111.9238, 55.98486, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643703, 5629877, 10.42881, 111.4609, 56.36318, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643759, 5629935, 10.41172, 110.8369, 55.82409, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643816, 5629991, 10.32814, 111.3351, 54.09827, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643872, 5630048, 10.36121, 110.9372, 53.59043, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _,
  1643927, 5630108, 10.38214, 111.1208, 54.36327, _ ;

 jsrc_noise =
  851.5497,
  1334.176,
  851.7628,
  1333.763,
  850.7783,
  1334.407,
  851.3549,
  1334.604,
  851.6039,
  1334.059,
  852.0295,
  1334.351,
  851.5128,
  1334.632,
  851.7574,
  1334.235,
  851.6926,
  1334.123,
  852.2081,
  1333.977,
  851.5474,
  1333.309,
  852.3996,
  1333.003,
  851.8854,
  1334.323,
  852.0712,
  1334.182,
  852.8131,
  1333.978,
  851.8556,
  1334.473,
  851.277,
  1334.323,
  851.7197,
  1333.239,
  851.713,
  1333.394,
  851.1327,
  1332.731,
  850.1468,
  1331.851,
  850.8623,
  1332.388,
  850.6614,
  1334.117,
  851.5204,
  1334.42,
  851.8162,
  1333.42,
  851.4053,
  1333.456,
  851.6202,
  1333.489,
  851.5677,
  1333.806,
  852.425,
  1332.986,
  851.3555,
  1333.457,
  851.9053,
  1333.692,
  852.9982,
  1334.12,
  852.447,
  1334.268,
  851.7476,
  1334.673,
  852.1924,
  1334.084,
  852.2639,
  1334.124,
  851.1191,
  1334.585,
  851.5846,
  1334.264,
  851.9114,
  1334.509,
  851.6002,
  1334.868,
  851.5359,
  1334.665,
  851.6472,
  1334.824,
  851.8442,
  1334.157,
  852.3253,
  1333.805,
  852.6849,
  1333.324,
  852.1635,
  1333.055,
  852.0715,
  1334.553,
  852.2643,
  1334.283,
  852.5503,
  1333.073,
  852.6456,
  1333,
  851.3979,
  1333.529,
  852.0196,
  1333.638,
  852.5549,
  1333.577,
  852.5194,
  1333.656,
  850.8351,
  1333.691,
  851.7248,
  1334.038,
  852.2759,
  1334.087,
  851.6208,
  1334.444,
  851.4178,
  1333.702,
  851.5169,
  1333.733,
  851.6017,
  1333.79,
  851.8281,
  1333.813,
  852.1267,
  1333.833,
  851.4827,
  1333.701,
  851.7807,
  1333.788,
  852.2953,
  1333.746,
  852.8468,
  1333.933,
  852.7632,
  1333.888,
  851.9421,
  1333.54,
  852.2387,
  1333.676,
  852.6745,
  1333.024,
  852.6483,
  1333.875,
  851.6016,
  1334.5,
  852.1445,
  1333.759,
  852.6953,
  1333.43,
  851.542,
  1333.604,
  851.3511,
  1333.831,
  851.9049,
  1333.792,
  852.4985,
  1333.804,
  851.8414,
  1334.428,
  851.7168,
  1334.567,
  851.6736,
  1333.705,
  851.9373,
  1333.523,
  851.9376,
  1333.678,
  851.4035,
  1334.328,
  851.5768,
  1333.936,
  851.6242,
  1334.079,
  852.0628,
  1333.395,
  852.476,
  1333.468,
  851.9061,
  1334.202,
  852.3094,
  1334.549,
  852.3283,
  1333.931,
  852.8773,
  1333.266,
  852.5342,
  1334.155,
  852.0713,
  1334.067,
  852.5269,
  1333.906,
  853.0667,
  1333.413,
  852.0969,
  1333.182,
  851.5302,
  1333.597,
  851.9824,
  1333.517,
  852.4921,
  1333.238,
  852.1439,
  1333.654,
  851.2886,
  1334.336,
  852.0663,
  1334.466,
  852.29,
  1333.829,
  851.2794,
  1333.954,
  850.2858,
  1333.238,
  851.2414,
  1333.376,
  851.9474,
  1333.009,
  851.884,
  1332.969,
  851.0743,
  1333.865,
  850.7581,
  1332.666,
  851.3239,
  1333.595,
  851.699,
  1333.525,
  851.5251,
  1333.28,
  851.2835,
  1333.909,
  851.8604,
  1333.873,
  852.0001,
  1333.268,
  852.6165,
  1333.097,
  851.8604,
  1333.151,
  851.5886,
  1333.363,
  851.7534,
  1333.471,
  852.5248,
  1332.733,
  852.6897,
  1332.675,
  851.9888,
  1333.38,
  852.0652,
  1333.658,
  852.4432,
  1333.392,
  852.5782,
  1333.402,
  851.8558,
  1334.152,
  851.8359,
  1334.196,
  852.3427,
  1333.713,
  852.6059,
  1332.679,
  851.4338,
  1333.287,
  851.5585,
  1334.157,
  851.7852,
  1333.009,
  852.7489,
  1333.331,
  852.0795,
  1334.066,
  851.1039,
  1333.816,
  851.7707,
  1333.904,
  852.5911,
  1333.7,
  851.7953,
  1334.108,
  851.4171,
  1334.386,
  851.6165,
  1333.918,
  851.9572,
  1333.581,
  850.9366,
  1333.806,
  850.8959,
  1333.819,
  851.3425,
  1333.727,
  851.5311,
  1333.24,
  852.0074,
  1332.969,
  851.8005,
  1333.347,
  851.2159,
  1333.208,
  851.9484,
  1333.802,
  852.1081,
  1333.939,
  852.5615,
  1334.003,
  851.9926,
  1333.613,
  851.4056,
  1333.601,
  852.1622,
  1333.292,
  852.6049,
  1333.268,
  852.8779,
  1333.183,
  852.0281,
  1333.755,
  852.0283,
  1333.986,
  852.3099,
  1333.224,
  852.9721,
  1333.387,
  852.0107,
  1333.946,
  851.6138,
  1333.612,
  851.7869,
  1332.771,
  852.4282,
  1332.972,
  851.5849,
  1333.74,
  851.3332,
  1334.225,
  851.9309,
  1333.168,
  852.5082,
  1333.198,
  851.2383,
  1333.366,
  851.4672,
  1334.076,
  851.7676,
  1333.335,
  852.0742,
  1333.672,
  851.407,
  1334.648,
  851.2115,
  1334.278,
  851.6981,
  1334.298,
  852.153,
  1333.626,
  852.2222,
  1333.829,
  850.9917,
  1334.007,
  851.1597,
  1333.674,
  851.6719,
  1333.273,
  852.0623,
  1333.617,
  851.605,
  1334.177,
  851.1852,
  1334.144,
  851.7872,
  1333.526,
  852.2977,
  1333.406,
  852.2408,
  1333.261,
  851.6871,
  1334.018,
  851.3952,
  1334.114,
  852.1069,
  1333.951,
  852.6785,
  1333.392,
  852.5118,
  1334.194,
  851.6865,
  1334.318,
  851.6381,
  1333.26,
  852.2893,
  1333.281,
  852.2809,
  1333.151,
  852.6695,
  1333.619,
  851.9109,
  1333.672,
  852.0106,
  1333.158,
  852.6472,
  1332.949,
  853.0255,
  1333.491,
  851.877,
  1334.154,
  852.4498,
  1333.791,
  852.6179,
  1333.253,
  852.8058,
  1333.65,
  851.7786,
  1334.064,
  851.6938,
  1333.955,
  851.9334,
  1333.511,
  852.4033,
  1333.061,
  850.5536,
  1332.839,
  850.6955,
  1332.58,
  851.3956,
  1332.426,
  852.4336,
  1333.734,
  851.2337,
  1334.54,
  851.9149,
  1334.505,
  852.1384,
  1334.092,
  851.2134,
  1331.698,
  850.5117,
  1332.724,
  851.0878,
  1333.646,
  851.0742,
  1332.476,
  851.435,
  1331.762,
  851.9213,
  1333.158,
  851.3976,
  1334.448,
  851.6369,
  1333.902,
  851.4257,
  1332.621,
  851.048,
  1331.617,
  850.4487,
  1331.618,
  850.5449,
  1332.828,
  851.4195,
  1333.225,
  852.0104,
  1333.377,
  852.0234,
  1333.806,
  851.2239,
  1333.723,
  851.3857,
  1332.535,
  852.0268,
  1332.709,
  851.6884,
  1332.044,
  851.4749,
  1333.288,
  851.5435,
  1333.118,
  851.942,
  1333.513,
  852.2932,
  1333.15,
  852.4493,
  1333.866,
  852.1677,
  1334.006,
  851.9882,
  1333.736,
  852.1757,
  1333.391,
  851.9545,
  1332.254,
  851.0631,
  1332.935,
  851.0143,
  1333.151,
  851.7201,
  1333.435,
  852.5787,
  1333.554,
  852.9131,
  1333.638,
  851.4594,
  1333.34,
  851.7991,
  1333.229,
  851.954,
  1332.742,
  852.1061,
  1332.402,
  851.8633,
  1334.635,
  851.4067,
  1333.633,
  851.9152,
  1333.162,
  852.4062,
  1333.455,
  850.9556,
  1333.546,
  851.1171,
  1333.792,
  852.205,
  1334.102,
  852.8145,
  1334.384,
  852.0862,
  1334.488,
  850.9319,
  1333.814,
  850.9888,
  1332.499,
  852.0356,
  1332.992,
  851.7101,
  1334.147,
  851.485,
  1334.173,
  851.8638,
  1333.884,
  851.778,
  1333.458,
  851.9166,
  1333.93,
  851.4718,
  1334.465,
  851.6027,
  1334.693,
  851.4721,
  1333.774,
  852.4203,
  1333.409,
  851.547,
  1334.342,
  851.6064,
  1334.6,
  852.2032,
  1333.349,
  852.0383,
  1332.961,
  852.6186,
  1333.843,
  851.8724,
  1334.049,
  851.701,
  1334.122,
  852.0712,
  1333.534,
  852.5389,
  1333.596,
  852.1265,
  1333.442,
  851.7627,
  1333.527,
  851.6763,
  1333.593,
  852.0119,
  1333.438,
  852.2369,
  1332.86,
  852.5193,
  1334.273,
  851.9229,
  1333.975,
  852.108,
  1333.771,
  852.3723,
  1333.63,
  852.3516,
  1333.84,
  851.9553,
  1334.098,
  851.8051,
  1333.563,
  852.6718,
  1333.983,
  852.5692,
  1333.211,
  851.8157,
  1334.455,
  851.5619,
  1334.044,
  852.3262,
  1333.919,
  852.7068,
  1333.23,
  852.126,
  1334.134,
  851.8212,
  1334.683,
  852.5853,
  1334.516,
  852.1899,
  1333.129,
  851.3905,
  1333.859,
  851.362,
  1334.362,
  851.9443,
  1334.132,
  852.599,
  1334.072,
  851.8901,
  1334.418,
  851.3845,
  1334.638,
  851.9304,
  1334.697,
  851.9725,
  1333.719,
  851.6259,
  1333.222,
  851.0075,
  1333.905,
  851.7493,
  1334.625,
  519.7802,
  -64.28521,
  519.6546,
  -64.66864,
  519.6701,
  -63.41517,
  519.8539,
  -63.842,
  519.6025,
  -64.48195,
  519.8022,
  -64.73811,
  519.8862,
  -64.03316,
  519.8618,
  -64.53721,
  519.7672,
  -64.30668,
  519.8412,
  -64.98522,
  519.2916,
  -64.62182,
  519.3942,
  -65.30912,
  519.8595,
  -64.54221,
  519.8901,
  -64.71459,
  519.8154,
  -65.41842,
  519.8392,
  -64.34736,
  519.675,
  -64.07482,
  519.5275,
  -64.80467,
  519.3763,
  -64.80488,
  519.2479,
  -64.59169,
  518.5397,
  -64.40399,
  518.9365,
  -64.56287,
  519.4427,
  -63.76083,
  519.6937,
  -64.30432,
  519.3564,
  -64.86456,
  519.4211,
  -64.86903,
  519.5379,
  -64.78953,
  519.5488,
  -64.54357,
  519.434,
  -65.70343,
  519.5198,
  -64.1963,
  519.634,
  -64.89812,
  519.8252,
  -65.51267,
  519.8546,
  -64.91907,
  519.8517,
  -64.17598,
  519.907,
  -64.91131,
  519.6384,
  -64.86545,
  519.6287,
  -63.7171,
  519.7628,
  -64.13966,
  519.8553,
  -64.38509,
  519.8579,
  -63.88451,
  519.8165,
  -63.92456,
  520.0143,
  -64.00154,
  519.7037,
  -64.53625,
  519.6889,
  -64.9436,
  519.6561,
  -65.43903,
  519.4431,
  -65.15311,
  519.7784,
  -64.55721,
  519.8908,
  -64.79597,
  519.5911,
  -65.71061,
  519.4147,
  -65.53185,
  519.4458,
  -64.02268,
  519.5652,
  -64.86841,
  519.6648,
  -65.42633,
  519.5977,
  -65.20053,
  519.5623,
  -63.65678,
  519.8153,
  -64.30057,
  519.8165,
  -64.87191,
  519.723,
  -64.06203,
  519.6648,
  -64.4756,
  519.5314,
  -64.41013,
  519.6109,
  -64.47796,
  519.7434,
  -64.61076,
  519.7136,
  -64.99113,
  519.6154,
  -64.2502,
  519.6818,
  -64.62143,
  519.8068,
  -64.91441,
  519.8793,
  -65.30537,
  519.8202,
  -65.13473,
  519.5635,
  -64.52541,
  519.5995,
  -65.04187,
  519.4946,
  -65.73891,
  519.6456,
  -65.27362,
  519.7908,
  -64.13757,
  519.5517,
  -64.91679,
  519.7275,
  -65.46037,
  519.5765,
  -64.34696,
  519.535,
  -64.03576,
  519.8119,
  -64.70412,
  519.6951,
  -65.16233,
  519.739,
  -64.52135,
  519.7821,
  -64.10966,
  519.6428,
  -64.54873,
  519.6032,
  -64.95603,
  519.6224,
  -64.95654,
  519.6882,
  -63.99006,
  519.5891,
  -64.34233,
  519.4331,
  -64.41148,
  519.3677,
  -65.18776,
  519.5643,
  -65.22095,
  519.7322,
  -64.44492,
  519.9083,
  -64.76956,
  519.8033,
  -64.99768,
  519.7544,
  -65.74144,
  519.7823,
  -65.10925,
  519.7333,
  -64.73656,
  519.7772,
  -65.14008,
  519.7048,
  -65.9931,
  519.4538,
  -65.12003,
  519.5204,
  -64.42334,
  519.7379,
  -64.70975,
  519.6737,
  -65.48908,
  519.6423,
  -64.99223,
  519.5602,
  -64.14556,
  519.5836,
  -64.88762,
  519.7009,
  -65.29745,
  519.5546,
  -64.31815,
  519.3743,
  -63.71979,
  519.4335,
  -64.61935,
  519.2815,
  -65.15148,
  519.2932,
  -64.81239,
  519.3652,
  -64.08134,
  519.0314,
  -64.37772,
  519.2619,
  -64.75968,
  519.4149,
  -64.99511,
  519.3351,
  -64.87889,
  519.5189,
  -64.1451,
  519.6989,
  -64.74201,
  519.6334,
  -65.23111,
  519.2404,
  -65.76547,
  519.4161,
  -64.97382,
  519.5562,
  -64.66821,
  519.3792,
  -64.61378,
  519.3951,
  -65.78966,
  519.4492,
  -65.98011,
  519.4615,
  -65.27163,
  519.6588,
  -65.08557,
  519.5052,
  -65.46244,
  519.5891,
  -65.69721,
  519.6517,
  -64.4816,
  519.8487,
  -64.6898,
  519.717,
  -65.25816,
  519.5002,
  -65.76576,
  519.2051,
  -64.50723,
  519.6624,
  -64.33996,
  519.3002,
  -64.79549,
  519.5312,
  -65.61179,
  519.6697,
  -64.73849,
  519.3495,
  -63.97675,
  519.4888,
  -64.71867,
  519.6259,
  -65.24891,
  519.6483,
  -64.38308,
  519.8994,
  -64.19482,
  519.7873,
  -64.34406,
  519.5423,
  -64.9282,
  519.4064,
  -63.93113,
  519.3761,
  -63.90613,
  519.4441,
  -64.14398,
  519.5666,
  -64.87122,
  519.4445,
  -65.15163,
  519.6024,
  -64.61747,
  519.2726,
  -64.36635,
  519.5041,
  -64.92031,
  519.5461,
  -65.31551,
  519.8532,
  -65.47117,
  519.5615,
  -64.65985,
  519.3996,
  -64.47256,
  519.4205,
  -64.98801,
  519.386,
  -65.72988,
  519.4802,
  -66.21149,
  519.6744,
  -64.94713,
  519.6096,
  -64.84073,
  519.4857,
  -65.4603,
  519.4763,
  -65.991,
  519.4877,
  -64.71246,
  519.4479,
  -64.56097,
  519.207,
  -65.15979,
  519.4111,
  -65.72861,
  519.4402,
  -64.48747,
  519.663,
  -64.41446,
  519.5642,
  -65.148,
  519.4908,
  -65.61143,
  519.1857,
  -64.71532,
  519.521,
  -64.30328,
  519.5034,
  -64.69628,
  519.6464,
  -65.21543,
  519.91,
  -63.85099,
  519.6807,
  -63.81718,
  519.7567,
  -64.49311,
  519.5383,
  -65.00141,
  519.5974,
  -64.90575,
  519.378,
  -63.86211,
  519.3093,
  -63.94358,
  519.2316,
  -64.95712,
  519.6579,
  -65.31467,
  519.7494,
  -64.57188,
  519.6158,
  -64.15247,
  519.4277,
  -64.83072,
  519.3632,
  -65.40605,
  519.2557,
  -65.14503,
  519.6674,
  -64.59401,
  519.6108,
  -64.49847,
  519.683,
  -65.08818,
  519.7249,
  -65.38684,
  519.6995,
  -65.18202,
  519.8093,
  -64.29969,
  519.6298,
  -64.72351,
  519.6848,
  -65.15885,
  519.4795,
  -65.1748,
  519.6439,
  -65.33092,
  519.4922,
  -64.7554,
  519.3016,
  -65.36372,
  519.4746,
  -65.64501,
  519.7414,
  -65.74952,
  519.6988,
  -64.49063,
  519.7921,
  -65.09763,
  519.5648,
  -65.42919,
  519.5931,
  -65.56893,
  519.6761,
  -64.3959,
  519.6067,
  -64.58701,
  519.4716,
  -65.10822,
  519.1008,
  -65.58367,
  518.9952,
  -64.04258,
  519.1182,
  -64.5162,
  519.127,
  -65.03859,
  519.5718,
  -65.30177,
  519.6617,
  -63.89734,
  519.633,
  -64.23932,
  519.5454,
  -64.84467,
  518.8149,
  -65.35345,
  519.0786,
  -63.99197,
  519.4317,
  -64.11294,
  519.1652,
  -64.47636,
  519.0493,
  -65.16273,
  519.4692,
  -65.31672,
  519.579,
  -64.12459,
  519.5222,
  -64.52475,
  518.9025,
  -64.87633,
  519.0333,
  -65.13192,
  518.6634,
  -64.87079,
  518.9929,
  -64.06666,
  519.0051,
  -64.72387,
  519.2665,
  -64.99319,
  519.5461,
  -64.87727,
  519.52,
  -64.28239,
  519.1118,
  -64.96161,
  519.0757,
  -65.18427,
  519.011,
  -65.40358,
  519.407,
  -64.8838,
  519.2115,
  -64.74119,
  519.497,
  -65.01114,
  519.5109,
  -65.37376,
  519.8886,
  -65.07843,
  519.8279,
  -64.84489,
  519.5349,
  -64.77406,
  519.3699,
  -65.33438,
  518.9561,
  -65.80765,
  518.9268,
  -64.687,
  519.168,
  -64.3685,
  519.4934,
  -64.95905,
  519.639,
  -65.56664,
  519.5311,
  -65.76082,
  519.1941,
  -64.63395,
  519.3852,
  -64.66651,
  519.1432,
  -65.26411,
  518.8606,
  -65.69324,
  519.7087,
  -64.44773,
  519.5456,
  -64.4073,
  519.4763,
  -65.04738,
  519.6891,
  -65.4501,
  519.2885,
  -63.92937,
  519.4232,
  -64.08545,
  519.6456,
  -64.83118,
  519.7874,
  -65.26269,
  519.6841,
  -64.6958,
  519.3282,
  -63.99442,
  518.864,
  -64.48833,
  519.4149,
  -65.18848,
  519.623,
  -64.66851,
  519.769,
  -64.26911,
  519.7789,
  -64.78822,
  519.4631,
  -64.87582,
  519.556,
  -64.79758,
  519.4897,
  -64.09717,
  519.778,
  -63.99515,
  519.48,
  -64.45,
  519.4949,
  -65.3895,
  519.6622,
  -64.18909,
  519.9698,
  -64.13309,
  519.5684,
  -65.05582,
  519.1638,
  -65.16589,
  519.7028,
  -65.28419,
  519.597,
  -64.6824,
  519.8127,
  -64.30213,
  519.5604,
  -64.8028,
  519.7018,
  -65.30223,
  519.4879,
  -65.40703,
  519.3834,
  -65.04025,
  519.4743,
  -64.65274,
  519.5764,
  -65.34512,
  519.3295,
  -65.91901,
  519.931,
  -65.35584,
  519.7925,
  -64.8234,
  519.6993,
  -64.90598,
  519.7782,
  -65.36382,
  519.7933,
  -65.18515,
  519.8298,
  -64.79614,
  519.5497,
  -64.65611,
  519.7551,
  -65.35136,
  519.5038,
  -65.7621,
  519.8785,
  -64.56815,
  519.6054,
  -64.59915,
  519.7165,
  -64.9603,
  519.6195,
  -65.65733,
  519.7383,
  -64.65781,
  519.8711,
  -64.176,
  519.8923,
  -64.81945,
  519.5141,
  -65.32977,
  519.65,
  -64.28492,
  519.8008,
  -63.96609,
  519.7262,
  -64.51041,
  519.8004,
  -65.1963,
  519.7828,
  -64.50761,
  519.7635,
  -63.89323,
  519.8181,
  -64.45503,
  519.5321,
  -64.99551,
  519.35,
  -64.98746,
  519.5178,
  -63.89922,
  519.8635,
  -64.16969,
  97.78869,
  -296.2242,
  97.32874,
  -296.189,
  98.38185,
  -295.6939,
  98.15433,
  -296.0852,
  97.58721,
  -296.2755,
  97.45293,
  -296.4019,
  98.12043,
  -296.0403,
  97.63965,
  -296.1761,
  97.8474,
  -296.2304,
  97.23103,
  -296.4817,
  97.20521,
  -296.3142,
  96.66426,
  -296.4922,
  97.64149,
  -296.2845,
  97.561,
  -296.3621,
  96.79958,
  -296.5909,
  97.76905,
  -296.1624,
  98.05083,
  -295.9063,
  97.3813,
  -296.1327,
  97.12123,
  -296.1629,
  97.49383,
  -296.0043,
  97.76391,
  -295.54,
  97.47395,
  -295.7597,
  98.33752,
  -295.7967,
  97.64616,
  -296.1936,
  97.29415,
  -296.1773,
  97.52258,
  -296.2489,
  97.32834,
  -296.2009,
  97.53976,
  -295.9153,
  96.69438,
  -296.601,
  97.69356,
  -296.1923,
  97.36287,
  -296.2824,
  96.77269,
  -296.7282,
  97.28857,
  -296.4164,
  98.04126,
  -296.1071,
  97.46051,
  -296.3786,
  97.36913,
  -296.1954,
  98.26553,
  -295.5973,
  98.00439,
  -296.0436,
  97.85672,
  -296.1787,
  98.1736,
  -295.9427,
  98.2467,
  -295.9775,
  98.25191,
  -295.9647,
  97.86069,
  -296.1624,
  97.22234,
  -296.3065,
  96.79589,
  -296.4549,
  97.05755,
  -296.2964,
  97.75378,
  -296.1591,
  97.54385,
  -296.4293,
  96.72215,
  -296.6262,
  96.59352,
  -296.5553,
  97.89097,
  -295.6678,
  97.46032,
  -296.1545,
  96.95181,
  -296.4969,
  96.97573,
  -296.4148,
  98.31319,
  -295.7444,
  97.85769,
  -296.1917,
  97.29788,
  -296.3519,
  98.16043,
  -295.8747,
  97.71295,
  -295.9031,
  97.78703,
  -296.0421,
  97.70956,
  -296.1366,
  97.41636,
  -296.2334,
  97.15981,
  -296.4283,
  97.7081,
  -295.8509,
  97.59474,
  -296.1248,
  97.34794,
  -296.389,
  97.02536,
  -296.5974,
  97.05659,
  -296.5301,
  97.37784,
  -296.1984,
  97.18707,
  -296.4121,
  96.63385,
  -296.6116,
  97.01777,
  -296.5601,
  98.09141,
  -296.124,
  97.38354,
  -296.2957,
  96.76901,
  -296.6136,
  97.75146,
  -295.9933,
  98.05903,
  -295.8178,
  97.27544,
  -296.2375,
  97.05018,
  -296.4036,
  97.89421,
  -296.0703,
  98.05622,
  -295.8625,
  97.71998,
  -296.1046,
  97.31636,
  -296.2448,
  97.38177,
  -296.0984,
  98.11709,
  -295.781,
  97.91559,
  -295.9578,
  97.82832,
  -296.0008,
  96.89853,
  -296.3491,
  96.97137,
  -296.3645,
  97.74601,
  -296.1007,
  97.58506,
  -296.2989,
  97.36658,
  -296.3735,
  96.63857,
  -296.7162,
  97.21918,
  -296.3956,
  97.61425,
  -296.2461,
  97.08059,
  -296.4693,
  96.48267,
  -296.786,
  97.20245,
  -296.4005,
  97.75945,
  -295.9477,
  97.44152,
  -296.1701,
  96.75069,
  -296.5128,
  97.06865,
  -296.2719,
  97.93751,
  -295.7009,
  97.52421,
  -296.1108,
  97.05876,
  -296.3203,
  97.92332,
  -295.6617,
  98.29586,
  -295.5572,
  97.52566,
  -296.0786,
  97.03057,
  -296.3272,
  97.22793,
  -296.0028,
  98.0322,
  -295.481,
  97.80647,
  -295.6678,
  97.6408,
  -295.7863,
  97.24112,
  -296.3152,
  97.14822,
  -296.0674,
  97.95609,
  -295.8737,
  97.57742,
  -296.2065,
  97.1929,
  -296.5404,
  96.63118,
  -296.616,
  97.22211,
  -296.1705,
  97.52509,
  -295.9342,
  97.35456,
  -295.9013,
  96.46004,
  -296.5614,
  96.06716,
  -296.7097,
  97.10645,
  -296.1999,
  97.35378,
  -296.1528,
  97.02036,
  -296.4702,
  96.73281,
  -296.4454,
  97.7626,
  -295.9407,
  97.68365,
  -296.1871,
  97.16684,
  -296.35,
  96.58839,
  -296.5199,
  97.44777,
  -295.8601,
  97.89383,
  -295.9692,
  97.34893,
  -295.8603,
  96.77998,
  -296.4373,
  97.46515,
  -296.0812,
  98.02604,
  -295.855,
  97.63116,
  -296.0759,
  96.96819,
  -296.3794,
  97.7562,
  -295.9253,
  98.05122,
  -295.9433,
  97.88132,
  -296.0829,
  97.33701,
  -296.1543,
  98.09096,
  -295.7138,
  98.37474,
  -295.6791,
  97.80466,
  -295.8145,
  97.38881,
  -295.8855,
  96.94583,
  -296.2391,
  97.43784,
  -295.9374,
  97.92736,
  -295.7077,
  97.54253,
  -296.0428,
  97.15142,
  -296.2413,
  97.04242,
  -296.5592,
  97.51492,
  -296.1449,
  97.87137,
  -295.8214,
  97.12134,
  -296.1765,
  96.77264,
  -296.5127,
  96.27258,
  -296.8915,
  97.27122,
  -296.3507,
  97.25357,
  -296.1627,
  96.96644,
  -296.318,
  96.35323,
  -296.6678,
  97.34989,
  -296.1579,
  97.47594,
  -296.0561,
  97.17244,
  -296.2006,
  96.59775,
  -296.5071,
  97.71026,
  -296.0652,
  97.99982,
  -295.7615,
  97.31155,
  -296.0033,
  96.79822,
  -296.5331,
  97.69839,
  -295.8829,
  97.84579,
  -295.7346,
  97.47203,
  -296.0498,
  97.28355,
  -296.1713,
  98.36678,
  -295.7506,
  98.2817,
  -295.6772,
  97.89639,
  -295.9938,
  97.2075,
  -296.2619,
  97.29594,
  -296.3711,
  98.338,
  -295.7036,
  97.97358,
  -295.4991,
  97.22012,
  -295.9013,
  96.79734,
  -296.4706,
  97.73474,
  -296.0563,
  97.94424,
  -295.6853,
  97.50318,
  -295.9117,
  96.96052,
  -296.4188,
  97.00439,
  -296.3031,
  97.66106,
  -295.9341,
  97.8169,
  -295.8142,
  97.14977,
  -296.3469,
  96.90929,
  -296.411,
  97.10127,
  -296.2833,
  97.82673,
  -295.9328,
  97.45603,
  -295.9498,
  97.01398,
  -296.4095,
  96.70923,
  -296.361,
  97.00425,
  -296.3985,
  97.46593,
  -296.1134,
  96.9705,
  -296.1484,
  96.5014,
  -296.4117,
  96.67751,
  -296.5492,
  97.7601,
  -295.9779,
  97.27563,
  -296.305,
  96.83874,
  -296.4366,
  96.7336,
  -296.592,
  97.74578,
  -295.889,
  97.53532,
  -295.9297,
  96.83316,
  -296.2943,
  96.36259,
  -296.543,
  97.82459,
  -295.5595,
  97.66631,
  -295.6704,
  97.01443,
  -296.0492,
  96.88815,
  -296.3658,
  98.21601,
  -295.7728,
  97.84743,
  -295.8235,
  97.49265,
  -296.182,
  96.90064,
  -296.0414,
  97.88149,
  -295.6014,
  98.0454,
  -295.4908,
  97.43337,
  -295.5543,
  97.0279,
  -295.963,
  97.08794,
  -296.0395,
  98.05678,
  -295.8142,
  97.71618,
  -296.0334,
  97.22964,
  -295.9255,
  97.01805,
  -295.8551,
  97.19071,
  -295.6167,
  97.75681,
  -295.5001,
  97.47328,
  -295.9464,
  97.15999,
  -296.1302,
  97.35798,
  -296.4061,
  97.72429,
  -295.6256,
  97.24415,
  -295.8925,
  97.03094,
  -296.1269,
  96.86119,
  -296.2278,
  97.34718,
  -296.0101,
  97.32163,
  -296.0671,
  97.31638,
  -296.2912,
  96.91081,
  -296.2622,
  97.33044,
  -296.303,
  97.54316,
  -296.2542,
  97.53467,
  -296.1557,
  96.93607,
  -296.3135,
  96.45867,
  -296.2083,
  97.24282,
  -295.7905,
  97.45887,
  -295.6709,
  97.17267,
  -296.1236,
  96.7204,
  -296.5245,
  96.55636,
  -296.5439,
  97.4826,
  -295.7147,
  97.53072,
  -296.0448,
  96.83765,
  -296.1774,
  96.29567,
  -296.2517,
  97.70084,
  -295.9308,
  97.77848,
  -295.9388,
  97.18681,
  -296.107,
  96.91164,
  -296.3659,
  98.05626,
  -295.5709,
  97.94788,
  -295.6319,
  97.12635,
  -296.1338,
  96.92491,
  -296.517,
  97.48251,
  -296.073,
  97.98521,
  -295.615,
  97.4288,
  -295.7115,
  97.02055,
  -296.1152,
  97.78353,
  -295.864,
  98.02917,
  -295.9082,
  97.60637,
  -296.2098,
  97.39066,
  -296.0716,
  97.53774,
  -296.1299,
  98.32913,
  -295.7413,
  98.21963,
  -295.7722,
  97.7472,
  -296.0104,
  96.93062,
  -296.3942,
  98.11864,
  -295.8645,
  98.04227,
  -296.0215,
  97.29257,
  -296.2806,
  97.0612,
  -296.3119,
  97.13141,
  -296.4107,
  97.71686,
  -296.0036,
  97.88005,
  -296.0022,
  97.63915,
  -296.061,
  96.98928,
  -296.2577,
  97.16733,
  -296.2228,
  97.29404,
  -296.1646,
  97.3277,
  -296.0378,
  97.11646,
  -296.2477,
  96.80464,
  -296.2905,
  97.10436,
  -296.4114,
  97.58086,
  -296.1209,
  97.41631,
  -296.2105,
  96.98595,
  -296.3861,
  97.10445,
  -296.3289,
  97.6022,
  -296.1227,
  97.60061,
  -296.1835,
  97.05012,
  -296.4809,
  96.76064,
  -296.4977,
  97.83485,
  -296.0731,
  97.81599,
  -295.8578,
  97.35137,
  -296.3195,
  96.69047,
  -296.5394,
  97.58719,
  -296.1728,
  97.96935,
  -296.0722,
  97.67069,
  -296.2474,
  97.07877,
  -296.2807,
  97.93981,
  -295.828,
  98.20421,
  -295.8502,
  97.65548,
  -296.0493,
  97.12508,
  -296.4438,
  97.78471,
  -296.129,
  98.15974,
  -295.8127,
  97.89939,
  -296.0409,
  97.28072,
  -296.2708,
  97.14658,
  -296.1388,
  98.13809,
  -295.6744,
  98.02993,
  -295.956,
  -159.5753,
  -151.056,
  -159.8442,
  -150.7696,
  -158.8566,
  -151.3106,
  -159.3669,
  -151.4404,
  -159.5549,
  -151.0313,
  -159.8745,
  -150.8103,
  -159.2631,
  -151.3515,
  -159.6363,
  -151.0944,
  -159.5449,
  -151.1807,
  -160.1561,
  -150.8403,
  -159.7189,
  -150.6569,
  -160.3537,
  -150.4522,
  -159.6545,
  -151.1141,
  -159.896,
  -151.1002,
  -160.4542,
  -150.487,
  -159.4793,
  -151.1906,
  -159.2237,
  -151.452,
  -159.7668,
  -150.9466,
  -159.838,
  -150.917,
  -159.8699,
  -151.1027,
  -159.1809,
  -151.1505,
  -159.4951,
  -150.6344,
  -158.9461,
  -151.5694,
  -159.5208,
  -151.1863,
  -159.8704,
  -150.8813,
  -159.6548,
  -150.9726,
  -159.7053,
  -150.9369,
  -159.5497,
  -150.9323,
  -160.5407,
  -150.5939,
  -159.7245,
  -151.0362,
  -159.8737,
  -150.9288,
  -160.5305,
  -150.5098,
  -159.9261,
  -150.837,
  -159.3611,
  -151.3785,
  -159.901,
  -150.983,
  -159.8345,
  -150.7394,
  -158.8983,
  -151.4934,
  -159.2633,
  -151.2564,
  -159.4779,
  -151.1526,
  -159.2392,
  -151.3902,
  -159.1556,
  -151.4754,
  -159.1915,
  -151.5301,
  -159.6111,
  -151.1187,
  -159.9961,
  -150.776,
  -160.3463,
  -150.4342,
  -160.1295,
  -150.5781,
  -159.6156,
  -151.2132,
  -159.8691,
  -151.029,
  -160.4629,
  -150.373,
  -160.4611,
  -150.3869,
  -159.2289,
  -151.0305,
  -159.8365,
  -150.8581,
  -160.3438,
  -150.6961,
  -160.1952,
  -150.5247,
  -158.8988,
  -151.2358,
  -159.5175,
  -151.1865,
  -159.9324,
  -150.8677,
  -159.2141,
  -151.304,
  -159.5501,
  -151.0616,
  -159.3909,
  -151.1672,
  -159.528,
  -151.1436,
  -159.6626,
  -151.0444,
  -159.9324,
  -150.8669,
  -159.2946,
  -151.1143,
  -159.7832,
  -151.0156,
  -159.9223,
  -150.903,
  -160.2597,
  -150.7274,
  -160.1858,
  -150.7638,
  -159.6952,
  -150.9668,
  -160.0445,
  -150.8033,
  -160.4398,
  -150.3577,
  -160.1655,
  -150.5947,
  -159.2763,
  -151.2916,
  -159.9689,
  -150.8063,
  -160.4188,
  -150.5492,
  -159.5071,
  -151.0965,
  -159.1609,
  -151.2144,
  -159.7818,
  -150.7789,
  -160.1528,
  -150.5648,
  -159.4523,
  -151.12,
  -159.3009,
  -151.3186,
  -159.4922,
  -150.9993,
  -159.7693,
  -150.8343,
  -159.7784,
  -150.8495,
  -159.0826,
  -151.3677,
  -159.3484,
  -151.3546,
  -159.395,
  -151.0711,
  -160.0476,
  -150.6091,
  -160.16,
  -150.5794,
  -159.4367,
  -151.1955,
  -159.6927,
  -151.1132,
  -159.9281,
  -150.7815,
  -160.6092,
  -150.4747,
  -160.0469,
  -150.835,
  -159.7333,
  -151.0829,
  -160.1181,
  -150.79,
  -160.6676,
  -150.4061,
  -159.7859,
  -150.6564,
  -159.2971,
  -151.0398,
  -159.7015,
  -150.8214,
  -160.353,
  -150.458,
  -159.7424,
  -150.7662,
  -159.0559,
  -151.3986,
  -159.8252,
  -150.9308,
  -160.1383,
  -150.5707,
  -159.2727,
  -151.1882,
  -158.9387,
  -151.6275,
  -159.5693,
  -151.1931,
  -159.9871,
  -150.5307,
  -159.8051,
  -150.7315,
  -159.1679,
  -151.3155,
  -159.3691,
  -150.9165,
  -159.5189,
  -150.9754,
  -159.7981,
  -150.7984,
  -159.6397,
  -150.7018,
  -159.3668,
  -151.2442,
  -159.6511,
  -151.1514,
  -160.0332,
  -150.7334,
  -160.4106,
  -150.3605,
  -159.922,
  -150.8571,
  -159.5162,
  -151.0934,
  -159.5098,
  -150.7048,
  -160.4108,
  -150.1807,
  -160.6167,
  -150.0302,
  -159.8973,
  -150.6145,
  -159.6547,
  -150.9578,
  -160.1127,
  -150.8024,
  -160.3997,
  -150.5377,
  -159.3497,
  -151.0634,
  -159.4946,
  -151.0689,
  -160.0249,
  -150.8109,
  -160.4917,
  -150.2919,
  -159.3925,
  -150.9324,
  -159.4914,
  -151.2206,
  -160.0259,
  -150.7128,
  -160.3956,
  -150.4727,
  -159.6155,
  -151.0434,
  -158.8752,
  -151.3251,
  -159.6758,
  -151.1552,
  -160.0811,
  -150.6997,
  -159.376,
  -151.1622,
  -159.1531,
  -151.3924,
  -159.4625,
  -151.11,
  -159.7772,
  -150.8064,
  -158.7505,
  -151.4796,
  -158.949,
  -151.3332,
  -159.3333,
  -151.2978,
  -159.615,
  -150.9082,
  -160.2664,
  -150.5059,
  -159.6982,
  -150.9117,
  -158.8774,
  -151.366,
  -159.771,
  -151.0866,
  -160.1737,
  -150.8866,
  -160.4034,
  -150.7858,
  -159.7424,
  -150.9705,
  -159.4066,
  -151.232,
  -159.8545,
  -150.7832,
  -160.576,
  -150.5956,
  -160.7211,
  -150.2613,
  -159.8564,
  -150.8338,
  -159.9333,
  -150.6796,
  -160.1923,
  -150.6686,
  -160.7532,
  -150.2539,
  -159.5755,
  -150.8806,
  -159.6148,
  -151.0584,
  -159.9585,
  -150.7668,
  -160.5218,
  -150.4454,
  -159.4046,
  -151.1711,
  -159.3498,
  -151.3922,
  -159.7742,
  -150.867,
  -160.342,
  -150.4261,
  -159.6405,
  -151.113,
  -159.1746,
  -151.277,
  -159.5016,
  -150.8441,
  -160.0134,
  -150.7788,
  -158.9107,
  -151.4305,
  -159.0125,
  -151.3852,
  -159.4636,
  -151.3605,
  -159.7801,
  -150.8222,
  -159.7618,
  -150.847,
  -158.8661,
  -151.3208,
  -159.1015,
  -151.1644,
  -159.7196,
  -150.8836,
  -160.1387,
  -150.8561,
  -159.5336,
  -151.2124,
  -159.1216,
  -151.144,
  -159.8014,
  -150.8593,
  -160.004,
  -150.7519,
  -160.0239,
  -150.6107,
  -159.3469,
  -151.0133,
  -159.2461,
  -151.3151,
  -159.8407,
  -150.7392,
  -160.1952,
  -150.6904,
  -159.9751,
  -150.7831,
  -159.2807,
  -151.3264,
  -159.3651,
  -150.9247,
  -159.9358,
  -150.7891,
  -160.1823,
  -150.4528,
  -160.1283,
  -150.7121,
  -159.5903,
  -151.0083,
  -160.0689,
  -150.4069,
  -160.5502,
  -150.4467,
  -160.3696,
  -150.526,
  -159.435,
  -151.2276,
  -159.9808,
  -150.9123,
  -160.3083,
  -150.5617,
  -160.4296,
  -150.6441,
  -159.3893,
  -151.0542,
  -159.5983,
  -151.002,
  -160.0293,
  -150.5303,
  -160.2553,
  -150.1543,
  -158.8923,
  -151.1263,
  -159.1369,
  -151.091,
  -159.8124,
  -150.6378,
  -160.0755,
  -150.6192,
  -158.9347,
  -151.428,
  -159.3941,
  -151.2222,
  -159.6356,
  -150.8062,
  -159.7092,
  -150.4977,
  -158.8931,
  -151.2256,
  -159.1867,
  -151.3311,
  -159.4607,
  -150.8288,
  -160.064,
  -150.7285,
  -159.9402,
  -150.561,
  -159.1169,
  -151.44,
  -159.4025,
  -151.0716,
  -159.8232,
  -150.5743,
  -159.7997,
  -150.3129,
  -159.5323,
  -150.5271,
  -159.259,
  -150.9978,
  -159.6483,
  -150.8994,
  -160.1189,
  -150.8542,
  -159.9604,
  -150.9245,
  -159.1408,
  -151.2771,
  -159.4399,
  -150.8048,
  -160.0106,
  -150.7139,
  -160.069,
  -150.3994,
  -159.4946,
  -150.9972,
  -159.7118,
  -150.8352,
  -159.9066,
  -150.8299,
  -160.2222,
  -150.4391,
  -159.9428,
  -150.7251,
  -159.7618,
  -151.0687,
  -159.6164,
  -150.9538,
  -160.0081,
  -150.4258,
  -160.3234,
  -150.1297,
  -159.5866,
  -150.7717,
  -159.3314,
  -150.7453,
  -159.904,
  -150.7627,
  -160.3278,
  -150.4672,
  -160.4876,
  -150.2093,
  -159.5134,
  -150.755,
  -159.7134,
  -150.8428,
  -160.237,
  -150.4857,
  -160.5107,
  -150.0064,
  -159.4239,
  -151.0585,
  -159.3766,
  -151.1173,
  -159.8709,
  -150.7911,
  -160.1535,
  -150.5901,
  -158.974,
  -151.1843,
  -159.0911,
  -151.2588,
  -159.9265,
  -150.8304,
  -160.2613,
  -150.6348,
  -159.623,
  -151.0415,
  -159.1621,
  -151.1248,
  -159.5452,
  -151.0539,
  -159.8356,
  -150.6929,
  -159.4138,
  -151.1252,
  -159.1651,
  -151.3237,
  -159.6304,
  -150.9727,
  -159.7144,
  -150.9159,
  -159.6232,
  -150.9683,
  -159.0288,
  -151.3217,
  -158.998,
  -151.4302,
  -159.4501,
  -151.0131,
  -160.0647,
  -150.5987,
  -159.1423,
  -151.3393,
  -159.2105,
  -151.3637,
  -159.9233,
  -150.6507,
  -159.8112,
  -150.5595,
  -160.1331,
  -150.728,
  -159.5463,
  -150.9965,
  -159.2473,
  -151.1902,
  -159.6563,
  -150.9076,
  -160.1887,
  -150.6232,
  -159.9769,
  -150.624,
  -159.6635,
  -150.8266,
  -159.6779,
  -151.006,
  -160.1221,
  -150.6633,
  -160.399,
  -150.4584,
  -160.091,
  -150.6491,
  -159.6495,
  -151.1001,
  -159.8651,
  -151.0924,
  -160.0594,
  -150.7236,
  -160.0002,
  -150.7605,
  -159.5056,
  -151.0237,
  -159.5864,
  -151.0447,
  -160.1853,
  -150.7485,
  -160.277,
  -150.4682,
  -159.565,
  -151.2099,
  -159.4134,
  -151.1357,
  -159.9271,
  -150.9354,
  -160.3671,
  -150.4943,
  -159.596,
  -150.9446,
  -159.3126,
  -151.2952,
  -159.7871,
  -150.9179,
  -159.986,
  -150.584,
  -159.2834,
  -151.0526,
  -159.0497,
  -151.5026,
  -159.472,
  -151.0029,
  -160.0851,
  -150.7533,
  -159.437,
  -151.271,
  -159.0852,
  -151.5798,
  -159.5884,
  -151.2727,
  -159.7547,
  -150.8745,
  -159.5541,
  -150.6815,
  -158.8684,
  -151.309,
  -159.2301,
  -151.3931,
  -156.3122,
  60.97182,
  -156.2296,
  61.60086,
  -156.204,
  60.21061,
  -156.317,
  60.64019,
  -156.1541,
  61.12182,
  -156.2485,
  61.38223,
  -156.2775,
  60.68825,
  -156.2997,
  61.08392,
  -156.4626,
  60.82326,
  -156.2463,
  61.5943,
  -155.9413,
  61.43772,
  -156.123,
  62.10432,
  -156.3216,
  61.10249,
  -156.396,
  61.25625,
  -156.2361,
  62.01009,
  -156.2448,
  60.8589,
  -156.3278,
  60.64494,
  -156.1657,
  61.3422,
  -155.9646,
  61.44635,
  -156.0641,
  61.0776,
  -155.7801,
  60.72212,
  -156.1137,
  61.14292,
  -156.2556,
  60.31506,
  -156.3004,
  60.95322,
  -156.2388,
  61.56037,
  -156.638,
  61.50607,
  -156.1777,
  61.6045,
  -156.2229,
  61.18901,
  -156.0494,
  61.84082,
  -156.3438,
  60.88774,
  -156.2688,
  61.55966,
  -156.1281,
  62.09147,
  -156.1815,
  61.44614,
  -156.4368,
  60.63417,
  -156.3748,
  61.33541,
  -156.1995,
  61.3068,
  -156.2738,
  60.18823,
  -156.2747,
  60.80523,
  -156.455,
  60.97504,
  -156.418,
  60.57426,
  -156.3904,
  60.48987,
  -156.4926,
  60.42589,
  -156.4752,
  60.86536,
  -156.0824,
  61.41297,
  -156.1433,
  61.895,
  -156.1274,
  61.62483,
  -156.3523,
  61.04505,
  -156.3379,
  61.32596,
  -156.1109,
  62.05192,
  -156.127,
  62.11165,
  -156.2081,
  60.72221,
  -156.2256,
  61.10239,
  -156.0993,
  61.79805,
  -156.3651,
  61.65931,
  -156.4466,
  60.40869,
  -156.4286,
  60.76149,
  -156.271,
  61.45647,
  -156.3233,
  60.64961,
  -156.3336,
  60.85413,
  -156.3981,
  60.83621,
  -156.3652,
  60.85213,
  -156.4741,
  61.13188,
  -156.2386,
  61.46095,
  -156.3449,
  60.80409,
  -156.2088,
  61.03249,
  -156.2039,
  61.43161,
  -156.279,
  61.85101,
  -156.2075,
  61.70988,
  -156.2173,
  61.38007,
  -156.1769,
  61.56014,
  -156.2914,
  62.26931,
  -156.2645,
  61.71023,
  -156.4683,
  60.76343,
  -156.2199,
  61.35083,
  -156.138,
  62.14041,
  -156.1281,
  60.94948,
  -156.2972,
  60.59846,
  -156.2643,
  61.14961,
  -156.3033,
  61.76156,
  -156.3022,
  60.82872,
  -156.2173,
  60.635,
  -156.3181,
  60.96868,
  -156.264,
  61.37223,
  -156.2745,
  61.12509,
  -156.3638,
  60.57541,
  -156.534,
  60.87111,
  -156.3183,
  60.85168,
  -156.1627,
  61.60418,
  -156.1301,
  61.76431,
  -156.3049,
  60.95821,
  -156.4053,
  61.19631,
  -156.6694,
  61.32633,
  -156.2725,
  62.23458,
  -156.2569,
  61.60439,
  -156.3606,
  61.18218,
  -156.2821,
  61.69334,
  -156.2231,
  62.31902,
  -156.0915,
  61.70776,
  -156.2842,
  60.82582,
  -156.4126,
  61.22937,
  -156.2322,
  61.92372,
  -155.9951,
  61.60791,
  -156.3463,
  60.69013,
  -156.4769,
  61.29008,
  -156.2659,
  61.87918,
  -156.2869,
  60.68668,
  -156.3794,
  60.44969,
  -156.2115,
  61.22919,
  -156.2639,
  61.68506,
  -156.0367,
  61.46889,
  -156.088,
  60.69756,
  -156.1989,
  60.93823,
  -156.0862,
  61.29526,
  -156.1468,
  61.52274,
  -156.1495,
  61.62093,
  -156.5563,
  60.65094,
  -156.4932,
  61.10424,
  -156.2184,
  61.89665,
  -156.2005,
  62.30777,
  -156.0207,
  61.40055,
  -156.2782,
  61.11736,
  -156.5152,
  61.26314,
  -156.3163,
  61.96194,
  -155.9395,
  62.38012,
  -156.0824,
  61.47819,
  -156.2175,
  61.37957,
  -156.1799,
  61.8296,
  -156.1254,
  62.03448,
  -156.2332,
  60.87391,
  -156.4449,
  61.05061,
  -156.3611,
  61.58053,
  -156.0133,
  62.29456,
  -156.1131,
  60.97142,
  -156.3442,
  60.85786,
  -156.2159,
  61.36815,
  -156.121,
  61.98035,
  -156.1904,
  61.12873,
  -156.3377,
  60.44817,
  -156.1447,
  61.05581,
  -156.1639,
  61.71321,
  -156.1713,
  60.85197,
  -156.346,
  60.56237,
  -156.3757,
  61.00425,
  -156.2418,
  61.37833,
  -156.2677,
  60.5645,
  -156.4814,
  60.38969,
  -156.3914,
  60.92184,
  -156.1887,
  61.35447,
  -156.2352,
  61.92103,
  -156.2355,
  61.1375,
  -156.4091,
  60.65068,
  -156.3253,
  61.37467,
  -156.0203,
  61.55311,
  -156.2401,
  61.66151,
  -156.2541,
  61.16217,
  -156.1755,
  60.79037,
  -156.2399,
  61.619,
  -156.1552,
  62.19656,
  -156.0897,
  62.48482,
  -156.4166,
  61.40149,
  -156.2775,
  61.32256,
  -156.109,
  61.93466,
  -156.2122,
  62.47007,
  -156.2192,
  61.43716,
  -156.2824,
  61.07066,
  -156.2692,
  61.62128,
  -156.1115,
  62.03065,
  -156.3342,
  61.06398,
  -156.4615,
  60.64377,
  -156.1465,
  61.51046,
  -156.3663,
  61.93159,
  -156.2309,
  60.75467,
  -156.2435,
  60.64568,
  -156.3887,
  61.19595,
  -156.2997,
  61.49468,
  -156.3319,
  60.3014,
  -156.2673,
  60.32854,
  -156.2816,
  60.90058,
  -156.2039,
  61.47077,
  -156.151,
  61.41646,
  -156.2354,
  60.09729,
  -156.3259,
  60.58216,
  -156.3019,
  61.33139,
  -156.1944,
  61.6343,
  -156.2817,
  60.83073,
  -156.3018,
  60.65822,
  -156.2444,
  61.29596,
  -156.283,
  61.81829,
  -156.2085,
  61.75756,
  -156.1054,
  61.11059,
  -156.2883,
  60.73642,
  -156.4905,
  61.21696,
  -156.22,
  61.79875,
  -156.1825,
  61.60145,
  -156.3149,
  60.96485,
  -156.2671,
  61.28434,
  -156.4542,
  61.62881,
  -155.9699,
  61.753,
  -156.1965,
  61.80108,
  -156.4046,
  61.00114,
  -156.2366,
  61.48104,
  -156.1427,
  62.12364,
  -156.3666,
  62.11037,
  -156.3599,
  60.9002,
  -156.3271,
  61.4615,
  -156.2895,
  61.93434,
  -156.1853,
  62.18913,
  -156.1513,
  60.84865,
  -156.2799,
  60.9063,
  -156.4671,
  61.85273,
  -156.1578,
  62.27953,
  -156.1683,
  60.85818,
  -156.14,
  60.989,
  -156.1002,
  61.66505,
  -156.0911,
  61.98956,
  -156.41,
  60.21362,
  -156.3469,
  60.7298,
  -156.508,
  61.27251,
  -156.0245,
  61.85633,
  -155.9647,
  60.61372,
  -156.0542,
  60.45575,
  -156.0313,
  60.72956,
  -156.1626,
  61.43996,
  -156.267,
  61.38025,
  -156.304,
  60.41305,
  -156.5337,
  60.81052,
  -156.1409,
  61.42868,
  -156.1771,
  61.80222,
  -155.8043,
  61.31782,
  -155.9919,
  60.86089,
  -156.2068,
  61.10007,
  -156.3362,
  61.75541,
  -156.1693,
  61.42267,
  -156.2035,
  60.70033,
  -156.0928,
  61.21303,
  -156.2142,
  61.37637,
  -156.0755,
  61.43955,
  -156.4524,
  61.32595,
  -156.4838,
  61.25901,
  -156.2845,
  61.52032,
  -156.0466,
  61.83622,
  -156.1601,
  61.30779,
  -156.3762,
  61.15352,
  -156.426,
  61.1028,
  -156.3849,
  61.59282,
  -155.9084,
  62.59351,
  -156.0287,
  61.56754,
  -156.1687,
  60.88136,
  -156.0026,
  61.52438,
  -156.1835,
  62.02795,
  -156.3012,
  62.25141,
  -156.265,
  60.9658,
  -156.3559,
  61.15923,
  -155.8962,
  61.70184,
  -155.9637,
  62.32875,
  -156.1478,
  60.94257,
  -156.2222,
  60.89307,
  -156.0937,
  61.4575,
  -156.0565,
  61.88727,
  -155.9588,
  60.42134,
  -156.1157,
  60.64515,
  -156.2126,
  61.34368,
  -156.3899,
  61.904,
  -156.3452,
  61.15543,
  -156.3162,
  60.64511,
  -156.085,
  61.00838,
  -156.1968,
  61.37259,
  -156.3166,
  61.01377,
  -156.325,
  60.59057,
  -156.311,
  61.19287,
  -156.1496,
  61.25079,
  -156.2888,
  61.13423,
  -156.2615,
  60.40107,
  -156.3503,
  60.61295,
  -156.2354,
  61.12474,
  -156.1422,
  61.75652,
  -156.1655,
  60.63294,
  -156.3454,
  60.55783,
  -156.2739,
  61.55257,
  -156.0377,
  61.70259,
  -156.2817,
  61.6818,
  -156.1323,
  61.01136,
  -156.2587,
  60.82043,
  -156.12,
  61.28264,
  -156.2292,
  61.75887,
  -156.1811,
  61.60903,
  -156.17,
  61.4217,
  -156.3202,
  61.20267,
  -156.2959,
  61.69818,
  -156.0684,
  62.03218,
  -156.2987,
  61.71641,
  -156.3264,
  61.16364,
  -156.3156,
  61.2961,
  -156.1386,
  61.69964,
  -156.1912,
  61.66279,
  -156.1746,
  61.07747,
  -156.2192,
  61.15613,
  -156.3277,
  61.73688,
  -156.2392,
  62.16626,
  -156.2009,
  61.0395,
  -156.2831,
  60.89991,
  -156.2838,
  61.47189,
  -156.1942,
  62.10273,
  -156.1962,
  61.08724,
  -156.322,
  60.67172,
  -156.4576,
  61.22912,
  -156.1799,
  61.78299,
  -156.1095,
  60.61647,
  -156.347,
  60.44319,
  -156.1804,
  61.04473,
  -156.2036,
  61.60485,
  -156.2803,
  60.91468,
  -156.2766,
  60.46131,
  -156.3233,
  60.86908,
  -156.4309,
  61.38142,
  -156.2627,
  61.35357,
  -156.1932,
  60.41601,
  -156.3184,
  60.76946,
  -9.135457,
  133.9586,
  -8.805316,
  134.0869,
  -9.868482,
  133.6278,
  -9.489536,
  133.8985,
  -8.987088,
  134.0178,
  -8.723711,
  134.1036,
  -9.53311,
  133.7651,
  -9.119905,
  134.0729,
  -9.249376,
  134.0144,
  -8.629782,
  134.2586,
  -8.746415,
  134.2146,
  -8.151993,
  134.3008,
  -9.120995,
  133.9065,
  -8.922902,
  134.1882,
  -8.187552,
  134.3051,
  -9.226713,
  133.7906,
  -9.532727,
  133.846,
  -8.831526,
  134.0662,
  -8.688764,
  134.0803,
  -8.897079,
  134.0356,
  -9.106925,
  133.5064,
  -8.881607,
  133.7197,
  -9.799979,
  133.4803,
  -9.430359,
  133.9336,
  -8.81442,
  134.0843,
  -9.136968,
  133.8725,
  -9.019121,
  134.0368,
  -8.989437,
  134.0301,
  -8.125579,
  134.2711,
  -9.31231,
  133.6934,
  -8.806966,
  134.0987,
  -8.16414,
  134.3985,
  -8.764901,
  134.0555,
  -9.420671,
  133.9322,
  -8.914673,
  134.0726,
  -8.80621,
  133.9488,
  -9.966488,
  133.5118,
  -9.423043,
  133.9164,
  -9.296165,
  134.0191,
  -9.609938,
  133.7022,
  -9.57583,
  133.6908,
  -9.719948,
  133.782,
  -9.242886,
  133.8711,
  -8.692471,
  134.153,
  -8.183899,
  134.3146,
  -8.592274,
  134.0943,
  -9.220564,
  133.9922,
  -8.919509,
  134.1958,
  -8.304423,
  134.3871,
  -8.048967,
  134.2889,
  -9.350272,
  133.7011,
  -9.119423,
  134.1027,
  -8.604239,
  134.327,
  -8.476886,
  134.1008,
  -9.737669,
  133.7802,
  -9.289804,
  134.0424,
  -8.674558,
  134.1097,
  -9.509874,
  133.7612,
  -9.287728,
  133.9099,
  -9.344876,
  133.8847,
  -9.188583,
  133.9424,
  -8.980599,
  134.0559,
  -8.621697,
  134.0865,
  -9.239202,
  133.718,
  -9.108131,
  134.106,
  -8.747596,
  134.0628,
  -8.423133,
  134.3206,
  -8.525249,
  134.2829,
  -8.794627,
  133.8771,
  -8.538258,
  134.2548,
  -7.94551,
  134.3924,
  -8.3967,
  134.118,
  -9.382429,
  133.8927,
  -8.805926,
  134.1851,
  -8.32414,
  134.3753,
  -9.237949,
  133.8132,
  -9.493939,
  133.7967,
  -8.96174,
  134.1397,
  -8.517042,
  134.202,
  -9.320601,
  133.8153,
  -9.520817,
  133.7101,
  -9.145827,
  134.0511,
  -8.707321,
  134.1405,
  -8.703221,
  133.9795,
  -9.565619,
  133.6192,
  -9.395402,
  133.8661,
  -9.297282,
  133.9849,
  -8.531776,
  134.1879,
  -8.415919,
  134.1359,
  -9.183751,
  133.9201,
  -9.068003,
  134.0555,
  -8.93585,
  134.2405,
  -8.149835,
  134.3895,
  -8.640676,
  134.1178,
  -9.015725,
  134.0403,
  -8.537457,
  134.1986,
  -7.922197,
  134.4862,
  -8.683231,
  134.0953,
  -9.250403,
  133.8663,
  -8.841889,
  134.259,
  -8.248546,
  134.357,
  -8.671762,
  134.0713,
  -9.638009,
  133.7552,
  -9.117782,
  134.1291,
  -8.411471,
  134.2338,
  -9.192921,
  133.8328,
  -9.622111,
  133.4262,
  -9.139234,
  133.8022,
  -8.655613,
  134.1857,
  -8.745235,
  134.0441,
  -9.439394,
  133.5657,
  -9.028032,
  133.7777,
  -9.009732,
  133.9739,
  -8.56612,
  134.3319,
  -8.729308,
  134.0637,
  -9.545493,
  133.7805,
  -9.050832,
  134.0832,
  -8.492682,
  134.1663,
  -8.019179,
  134.3495,
  -8.774204,
  134.0196,
  -9.231211,
  134.0382,
  -8.774663,
  134.0178,
  -8.239791,
  134.4015,
  -7.688596,
  134.5113,
  -8.584228,
  134.1628,
  -8.707961,
  134.1896,
  -8.36748,
  134.3663,
  -8.13982,
  134.3588,
  -9.253383,
  133.7684,
  -9.136901,
  133.953,
  -8.618269,
  134.2423,
  -8.036895,
  134.3363,
  -9.10666,
  133.8333,
  -9.434401,
  133.8918,
  -8.748071,
  134.0543,
  -8.169525,
  134.2176,
  -9.04096,
  133.8567,
  -9.500818,
  133.7192,
  -8.914635,
  134.0752,
  -8.446165,
  134.2067,
  -9.217649,
  133.7216,
  -9.604208,
  133.706,
  -9.213058,
  133.9634,
  -8.750359,
  134.0827,
  -9.624093,
  133.4111,
  -9.703143,
  133.5078,
  -9.290584,
  133.8951,
  -9.043874,
  134.0296,
  -8.434718,
  134.2433,
  -9.06848,
  133.8798,
  -9.43577,
  133.8673,
  -8.964247,
  134.0642,
  -8.725204,
  134.2351,
  -8.422403,
  134.285,
  -9.001907,
  134.0414,
  -9.360645,
  133.8673,
  -8.78661,
  134.223,
  -8.145827,
  134.4519,
  -7.854006,
  134.621,
  -8.880251,
  134.2251,
  -8.749851,
  134.2243,
  -8.379904,
  134.4341,
  -8.007271,
  134.4532,
  -8.75352,
  133.9758,
  -9.063841,
  134.0796,
  -8.699822,
  134.2651,
  -8.030319,
  134.5267,
  -9.119692,
  133.9533,
  -9.381047,
  133.9124,
  -8.660367,
  134.1346,
  -8.229873,
  134.3952,
  -9.079798,
  133.6186,
  -9.480832,
  133.7843,
  -9.15014,
  133.908,
  -8.851923,
  134.181,
  -9.822231,
  133.6669,
  -9.80636,
  133.6657,
  -9.290484,
  133.9888,
  -8.652536,
  134.2036,
  -8.849488,
  134.0677,
  -9.98547,
  133.6276,
  -9.586432,
  133.7449,
  -8.944204,
  134.0852,
  -8.589804,
  134.2414,
  -9.38482,
  133.8985,
  -9.58559,
  133.6772,
  -8.98273,
  134.0061,
  -8.62752,
  134.3836,
  -8.60228,
  134.1926,
  -9.204787,
  133.938,
  -9.433572,
  133.7772,
  -8.881431,
  134.2329,
  -8.421125,
  134.1541,
  -8.618167,
  134.0373,
  -9.319454,
  133.9572,
  -8.813386,
  134.0133,
  -8.61704,
  134.3141,
  -8.395185,
  134.1332,
  -8.524384,
  134.2043,
  -9.170566,
  134.0323,
  -8.494421,
  134.069,
  -8.029476,
  134.4852,
  -8.134211,
  134.4672,
  -9.234982,
  133.8789,
  -8.89842,
  134.1585,
  -8.421836,
  134.3355,
  -8.168087,
  134.3884,
  -9.271252,
  133.7272,
  -9.333386,
  134.068,
  -8.664001,
  134.4273,
  -8.31499,
  134.3351,
  -9.475629,
  133.6161,
  -9.310398,
  133.7096,
  -8.687313,
  134.1859,
  -8.403937,
  134.2155,
  -9.86432,
  133.495,
  -9.538321,
  133.7955,
  -8.953585,
  134.0355,
  -8.446996,
  133.8113,
  -9.52275,
  133.6306,
  -9.63502,
  133.5925,
  -9.348933,
  134.1577,
  -8.730947,
  134.2247,
  -8.669488,
  134.1016,
  -9.704088,
  133.7331,
  -9.410659,
  133.9537,
  -8.623412,
  134.2572,
  -8.444605,
  134.1271,
  -8.811094,
  133.763,
  -9.162573,
  133.7394,
  -8.961413,
  134.1673,
  -8.749318,
  134.1645,
  -8.719611,
  134.0016,
  -9.341789,
  133.4451,
  -8.602629,
  133.9833,
  -8.647351,
  134.0918,
  -8.632836,
  134.1416,
  -8.772613,
  133.9892,
  -8.884159,
  133.9324,
  -8.787015,
  134.0805,
  -8.26565,
  134.2715,
  -8.722037,
  134.1129,
  -9.033588,
  134.0336,
  -9.081685,
  134.1096,
  -8.587768,
  134.3165,
  -7.905381,
  134.356,
  -8.792418,
  134.0167,
  -9.213684,
  133.8614,
  -8.688154,
  134.0137,
  -8.170286,
  134.3549,
  -8.135158,
  134.3636,
  -9.013107,
  133.6998,
  -9.085229,
  134.0964,
  -8.516309,
  134.2346,
  -7.908556,
  134.3448,
  -9.196762,
  133.8674,
  -9.229192,
  133.9246,
  -8.657224,
  134,
  -8.331236,
  134.1113,
  -9.51639,
  133.5718,
  -9.4511,
  133.6728,
  -8.732771,
  134.2286,
  -8.327967,
  134.4118,
  -8.923436,
  134.0251,
  -9.329226,
  133.7502,
  -9.028307,
  133.7716,
  -8.651619,
  134.1431,
  -9.165346,
  133.8029,
  -9.500083,
  133.8171,
  -9.119481,
  133.919,
  -8.74646,
  133.9271,
  -8.971452,
  133.9798,
  -9.642523,
  133.6467,
  -9.589424,
  133.7241,
  -9.173183,
  133.8998,
  -8.535812,
  134.2532,
  -9.504222,
  133.7561,
  -9.586291,
  133.8208,
  -8.488228,
  134.222,
  -8.580844,
  134.0997,
  -8.590674,
  134.2617,
  -9.141512,
  133.8366,
  -9.356075,
  133.7722,
  -8.876314,
  134.0787,
  -8.407894,
  134.2198,
  -8.556447,
  134.182,
  -8.768678,
  134.1294,
  -8.829388,
  134.1365,
  -8.569503,
  134.1093,
  -8.234684,
  134.1499,
  -8.549394,
  134.2115,
  -9.016842,
  133.9851,
  -8.93368,
  134.0353,
  -8.564446,
  134.1878,
  -8.619871,
  134.1311,
  -9.153317,
  133.8945,
  -9.270854,
  134.0921,
  -8.567855,
  134.2359,
  -8.251354,
  134.3268,
  -9.296835,
  133.9954,
  -9.218262,
  133.8025,
  -8.737812,
  134.2041,
  -8.178126,
  134.3913,
  -9.071939,
  133.7959,
  -9.529107,
  133.7968,
  -8.988797,
  134.1348,
  -8.477416,
  134.184,
  -9.30624,
  133.6021,
  -9.641342,
  133.7528,
  -9.181249,
  133.9558,
  -8.547865,
  134.1965,
  -9.269751,
  133.9094,
  -9.673532,
  133.6676,
  -9.368781,
  133.9689,
  -8.836574,
  134.1464,
  -8.701526,
  134.1147,
  -9.659003,
  133.5422,
  -9.477873,
  133.8292,
  96.64702,
  53.87895,
  96.86759,
  53.49522,
  95.89323,
  54.24051,
  96.33448,
  54.07492,
  96.62151,
  53.81536,
  96.89398,
  53.61079,
  96.24081,
  54.03342,
  96.68494,
  53.74918,
  96.5957,
  53.95713,
  97.04021,
  53.5111,
  96.77229,
  53.5672,
  97.37828,
  53.17188,
  96.64265,
  53.73263,
  96.94239,
  53.7731,
  97.38539,
  53.15443,
  96.40351,
  53.77769,
  96.25876,
  54.09082,
  96.80212,
  53.66111,
  96.89024,
  53.61305,
  96.68158,
  53.67017,
  96.39964,
  53.66671,
  96.56874,
  53.63207,
  95.85379,
  54.24902,
  96.50029,
  53.94798,
  96.97716,
  53.65685,
  96.64461,
  53.65199,
  96.73436,
  53.66461,
  96.67326,
  53.77733,
  97.47145,
  53.05394,
  96.40496,
  53.78531,
  96.93838,
  53.57451,
  97.43801,
  53.12495,
  96.86504,
  53.48197,
  96.41129,
  54.09932,
  96.97918,
  53.71471,
  96.82043,
  53.53782,
  95.90616,
  54.21993,
  96.29984,
  54.02094,
  96.64525,
  53.96315,
  96.17373,
  54.10739,
  96.10209,
  54.18088,
  96.13503,
  54.31259,
  96.61012,
  53.91549,
  96.96096,
  53.48646,
  97.31561,
  53.29549,
  96.94523,
  53.39967,
  96.52754,
  53.79864,
  96.84631,
  53.71458,
  97.40519,
  53.14158,
  97.46025,
  53.02666,
  96.29221,
  53.92485,
  96.78786,
  53.74121,
  97.19317,
  53.39726,
  96.9986,
  53.27936,
  96.0433,
  54.22172,
  96.58417,
  54.00617,
  96.98634,
  53.46666,
  96.18569,
  54.04127,
  96.52941,
  54.01624,
  96.3892,
  53.95347,
  96.46783,
  53.94199,
  96.76102,
  53.7792,
  96.9633,
  53.53269,
  96.42342,
  53.83627,
  96.81702,
  53.87919,
  96.92994,
  53.55653,
  97.22815,
  53.33337,
  97.16255,
  53.41538,
  96.76286,
  53.56822,
  97.0338,
  53.44678,
  97.46325,
  53.00691,
  97.04155,
  53.32346,
  96.35104,
  54.06827,
  96.8895,
  53.55029,
  97.3614,
  53.1877,
  96.44482,
  53.87259,
  96.24481,
  54.16481,
  96.74383,
  53.70443,
  97.14436,
  53.38289,
  96.38004,
  53.88499,
  96.12524,
  54.04486,
  96.62965,
  53.87481,
  97.06286,
  53.51779,
  96.73282,
  53.6448,
  96.1634,
  54.06758,
  96.52522,
  54.10102,
  96.46204,
  53.95407,
  97.00536,
  53.27327,
  97.11042,
  53.20876,
  96.49603,
  53.82591,
  96.71442,
  53.75773,
  96.94669,
  53.66817,
  97.53753,
  53.16065,
  96.9827,
  53.47435,
  96.73061,
  53.84836,
  97.15321,
  53.44464,
  97.61956,
  53.07003,
  96.90255,
  53.39827,
  96.42461,
  53.867,
  96.89398,
  53.6498,
  97.37128,
  53.23698,
  96.79183,
  53.54873,
  96.18315,
  54.25331,
  96.86581,
  53.90277,
  97.20206,
  53.30682,
  96.2476,
  53.90206,
  95.86059,
  54.09067,
  96.46753,
  53.77734,
  97.02757,
  53.5422,
  96.8905,
  53.67448,
  96.17626,
  53.98367,
  96.35218,
  53.96997,
  96.92174,
  53.79911,
  97.00765,
  53.49791,
  96.76988,
  53.53966,
  96.20673,
  54.10315,
  96.68922,
  53.87238,
  97.11374,
  53.4243,
  97.49072,
  53.15843,
  96.73139,
  53.54971,
  96.47629,
  54.00195,
  96.79929,
  53.60886,
  97.42571,
  53.07729,
  97.61314,
  52.92944,
  97.00909,
  53.4777,
  96.85353,
  53.6856,
  97.24443,
  53.31521,
  97.38966,
  53.24944,
  96.34148,
  53.79144,
  96.52309,
  53.89057,
  97.0727,
  53.54334,
  97.48786,
  53.03484,
  96.34961,
  53.72533,
  96.35938,
  54.04153,
  96.68723,
  53.48436,
  97.25336,
  53.18615,
  96.51708,
  53.67507,
  96.21527,
  54.06978,
  96.7085,
  53.62507,
  97.14545,
  53.29823,
  96.45296,
  53.76919,
  96.13883,
  54.08789,
  96.57083,
  53.81747,
  96.94221,
  53.54913,
  96.13799,
  54.07966,
  95.91902,
  54.21062,
  96.41119,
  53.9468,
  96.78959,
  53.69254,
  97.20551,
  53.45646,
  96.54154,
  53.6801,
  96.36398,
  54.09034,
  96.79597,
  53.75066,
  97.03465,
  53.5748,
  97.2161,
  53.38077,
  96.67397,
  53.69977,
  96.41595,
  54.03843,
  97.00555,
  53.62552,
  97.45506,
  53.2143,
  97.80662,
  52.9592,
  96.88012,
  53.70704,
  96.86877,
  53.68002,
  97.37357,
  53.37928,
  97.60499,
  53.05499,
  96.72742,
  53.64057,
  96.59653,
  54.00798,
  97.02154,
  53.53953,
  97.42753,
  53.08992,
  96.55828,
  53.88212,
  96.36878,
  54.03875,
  96.90504,
  53.56651,
  97.30447,
  53.25599,
  96.48523,
  53.65827,
  96.17878,
  54.04278,
  96.68509,
  53.75077,
  96.822,
  53.58644,
  95.97007,
  54.20083,
  95.95235,
  54.27504,
  96.52716,
  54.03114,
  96.92245,
  53.56248,
  96.82761,
  53.57005,
  95.96375,
  54.34246,
  96.3055,
  54.10231,
  96.79205,
  53.65866,
  97.07183,
  53.46865,
  96.46325,
  53.9838,
  96.23161,
  54.01941,
  96.80875,
  53.70501,
  97.12026,
  53.37077,
  97.15701,
  53.33998,
  96.57227,
  53.82545,
  96.3409,
  53.96688,
  96.90331,
  53.5849,
  97.17285,
  53.35528,
  96.98007,
  53.35673,
  96.52791,
  54.00579,
  96.81792,
  53.72931,
  97.1073,
  53.50181,
  97.20132,
  53.34257,
  97.07552,
  53.34497,
  96.70374,
  53.74261,
  97.06309,
  53.36117,
  97.46898,
  53.08167,
  97.55083,
  53.12767,
  96.53133,
  53.89431,
  96.95039,
  53.67654,
  97.2975,
  53.31109,
  97.39589,
  53.15074,
  96.37026,
  53.83324,
  96.76374,
  53.85136,
  97.19781,
  53.47216,
  97.38287,
  53.01285,
  96.13593,
  53.87077,
  96.42819,
  54.01876,
  96.8403,
  53.59753,
  97.14975,
  53.26606,
  95.85133,
  54.272,
  96.28233,
  54.01039,
  96.76755,
  53.66652,
  97.09746,
  53.00725,
  96.06603,
  53.86991,
  96.10011,
  53.95955,
  96.56047,
  54.00035,
  96.97103,
  53.4963,
  96.92615,
  53.44019,
  96.08788,
  54.20059,
  96.55474,
  54.00429,
  96.87663,
  53.56397,
  96.91508,
  53.49185,
  96.69376,
  53.698,
  96.40902,
  53.91849,
  96.69714,
  53.76483,
  96.9705,
  53.55806,
  96.88783,
  53.5592,
  96.18266,
  53.81021,
  96.71789,
  53.59085,
  97.03117,
  53.46511,
  97.02351,
  53.4139,
  96.68382,
  53.48247,
  96.57716,
  53.58493,
  96.82219,
  53.59773,
  97.21136,
  53.25978,
  96.86754,
  53.55514,
  96.73705,
  53.76072,
  96.72008,
  53.81272,
  97.18199,
  53.54074,
  97.57582,
  53.03568,
  96.68771,
  53.43079,
  96.55422,
  53.7734,
  96.94307,
  53.48628,
  97.52943,
  53.18549,
  97.47403,
  53.23972,
  96.47316,
  53.72628,
  96.75262,
  53.79195,
  97.16876,
  53.29689,
  97.64797,
  52.91267,
  96.43231,
  53.81736,
  96.58899,
  53.90601,
  96.91089,
  53.41924,
  97.18123,
  53.21349,
  96.01588,
  53.84572,
  96.18841,
  53.98294,
  96.9398,
  53.56201,
  97.41837,
  53.3959,
  96.73146,
  53.77011,
  96.19893,
  54.05309,
  96.51569,
  53.70632,
  96.80228,
  53.51662,
  96.42987,
  53.71776,
  96.18985,
  54.02875,
  96.58229,
  53.82766,
  96.76733,
  53.59195,
  96.64936,
  53.71112,
  95.96453,
  54.10201,
  96.19262,
  54.06142,
  96.68972,
  53.83073,
  97.08865,
  53.41349,
  96.21506,
  54.04187,
  96.21871,
  54.09161,
  97.00854,
  53.35272,
  97.01295,
  53.34519,
  97.14678,
  53.41835,
  96.49732,
  53.69056,
  96.43167,
  53.97525,
  96.91331,
  53.62441,
  97.18999,
  53.36354,
  96.9203,
  53.4687,
  96.77972,
  53.54855,
  96.87666,
  53.59909,
  97.11201,
  53.4137,
  97.3637,
  53.1273,
  97.10474,
  53.41452,
  96.64366,
  53.7933,
  96.89482,
  53.71804,
  97.16553,
  53.38324,
  96.99638,
  53.44564,
  96.56923,
  53.69914,
  96.70252,
  53.97455,
  97.19132,
  53.4897,
  97.35705,
  53.13908,
  96.51,
  53.87242,
  96.49865,
  53.88786,
  96.92491,
  53.57679,
  97.39471,
  53.10952,
  96.53465,
  53.65542,
  96.28519,
  53.97191,
  96.77134,
  53.6995,
  97.13009,
  53.30853,
  96.24915,
  53.84383,
  96.13412,
  54.16755,
  96.64586,
  53.82019,
  97.08936,
  53.39629,
  96.4371,
  53.83921,
  95.99113,
  54.13032,
  96.53549,
  53.95083,
  96.90091,
  53.62335,
  96.81501,
  53.55672,
  95.97681,
  54.05401,
  96.26982,
  54.08004,
  75.51859,
  -54.08709,
  75.23147,
  -54.5355,
  75.3961,
  -53.29797,
  75.55688,
  -53.68099,
  75.3566,
  -54.16922,
  75.26958,
  -54.45105,
  75.4162,
  -53.70248,
  75.38531,
  -54.14769,
  75.52645,
  -53.97329,
  75.34688,
  -54.61319,
  75.23702,
  -54.47147,
  75.20194,
  -55.06744,
  75.36372,
  -54.13785,
  75.45895,
  -54.3775,
  75.20199,
  -55.05239,
  75.33098,
  -53.94096,
  75.4597,
  -53.67615,
  75.36191,
  -54.39209,
  75.16953,
  -54.46145,
  75.36732,
  -54.21752,
  75.38213,
  -53.81436,
  75.37733,
  -54.05695,
  75.51015,
  -53.27807,
  75.45236,
  -53.79033,
  75.41233,
  -54.46706,
  75.37808,
  -54.19176,
  75.39451,
  -54.33945,
  75.39181,
  -54.1788,
  75.21043,
  -55.0731,
  75.40028,
  -53.98528,
  75.33826,
  -54.54152,
  75.25341,
  -55.15313,
  75.26748,
  -54.50189,
  75.55816,
  -53.80283,
  75.42896,
  -54.3552,
  75.16218,
  -54.35055,
  75.51836,
  -53.24767,
  75.4175,
  -53.84812,
  75.55477,
  -54.16561,
  75.42219,
  -53.66631,
  75.54333,
  -53.46295,
  75.58223,
  -53.52993,
  75.49554,
  -53.94402,
  75.32068,
  -54.61244,
  75.22739,
  -54.98266,
  75.21947,
  -54.63861,
  75.41308,
  -54.04442,
  75.45478,
  -54.39002,
  75.27288,
  -55.04627,
  75.12544,
  -55.18523,
  75.32343,
  -53.80637,
  75.39137,
  -54.30791,
  75.38635,
  -54.82091,
  75.21485,
  -54.68422,
  75.56799,
  -53.4447,
  75.61134,
  -53.93412,
  75.2687,
  -54.47602,
  75.34281,
  -53.5691,
  75.4961,
  -53.82009,
  75.39876,
  -53.8718,
  75.44255,
  -54.09045,
  75.41682,
  -54.20765,
  75.25925,
  -54.52288,
  75.31283,
  -53.82047,
  75.53893,
  -54.13307,
  75.31055,
  -54.48671,
  75.26873,
  -54.86162,
  75.35027,
  -54.76934,
  75.38833,
  -54.34781,
  75.36046,
  -54.65005,
  75.21769,
  -55.18739,
  75.20079,
  -54.65434,
  75.52124,
  -53.78849,
  75.31606,
  -54.48901,
  75.19054,
  -55.03466,
  75.32172,
  -53.92942,
  75.42559,
  -53.61789,
  75.33719,
  -54.26687,
  75.31184,
  -54.72097,
  75.32565,
  -53.86648,
  75.34958,
  -53.54819,
  75.46464,
  -54.10466,
  75.37309,
  -54.57225,
  75.31036,
  -54.39969,
  75.398,
  -53.56993,
  75.52962,
  -53.83891,
  75.44175,
  -53.93009,
  75.22988,
  -54.75896,
  75.17886,
  -54.80185,
  75.43018,
  -53.98878,
  75.42763,
  -54.18171,
  75.45654,
  -54.48278,
  75.26601,
  -55.15636,
  75.34913,
  -54.569,
  75.46776,
  -54.19893,
  75.3456,
  -54.75824,
  75.26219,
  -55.2667,
  75.23088,
  -54.58926,
  75.41037,
  -53.88054,
  75.50363,
  -54.37549,
  75.33134,
  -54.99093,
  75.26569,
  -54.39549,
  75.55569,
  -53.57841,
  75.5463,
  -54.2833,
  75.25081,
  -54.89548,
  75.41616,
  -53.79699,
  75.45458,
  -53.53382,
  75.39362,
  -54.10411,
  75.33014,
  -54.58737,
  75.35191,
  -54.41789,
  75.41148,
  -53.51297,
  75.43633,
  -53.90536,
  75.46191,
  -54.22391,
  75.49309,
  -54.52798,
  75.20796,
  -54.40123,
  75.43697,
  -53.60555,
  75.52506,
  -54.13408,
  75.33442,
  -54.64255,
  75.13214,
  -55.10266,
  75.18999,
  -54.40135,
  75.43524,
  -53.96434,
  75.26932,
  -54.18369,
  75.21095,
  -55.11829,
  75.13557,
  -55.37659,
  75.2363,
  -54.49734,
  75.41742,
  -54.48114,
  75.28939,
  -54.89066,
  75.1829,
  -55.10565,
  75.24188,
  -53.90519,
  75.52155,
  -54.08765,
  75.38099,
  -54.68324,
  75.08833,
  -55.16176,
  75.1459,
  -53.908,
  75.53945,
  -53.85357,
  75.35417,
  -54.55063,
  75.12238,
  -55.02716,
  75.30126,
  -54.11128,
  75.50228,
  -53.62773,
  75.39213,
  -54.24347,
  75.28555,
  -54.78887,
  75.28171,
  -53.92458,
  75.43966,
  -53.57539,
  75.47146,
  -53.9573,
  75.3376,
  -54.44309,
  75.46003,
  -53.50657,
  75.53117,
  -53.32923,
  75.49357,
  -53.80397,
  75.43829,
  -54.30436,
  75.31378,
  -54.77874,
  75.24023,
  -54.13256,
  75.52933,
  -53.80793,
  75.47945,
  -54.37497,
  75.39733,
  -54.57701,
  75.32053,
  -54.77999,
  75.34427,
  -54.1715,
  75.57262,
  -53.81448,
  75.43783,
  -54.56,
  75.28275,
  -55.18037,
  75.23969,
  -55.55927,
  75.50911,
  -54.37379,
  75.41422,
  -54.41987,
  75.34859,
  -54.86227,
  75.16001,
  -55.3903,
  75.21913,
  -54.26826,
  75.53616,
  -54.10493,
  75.39699,
  -54.67525,
  75.1858,
  -55.14968,
  75.42086,
  -54.06858,
  75.59429,
  -53.76233,
  75.31252,
  -54.48466,
  75.28884,
  -55.01132,
  75.30601,
  -53.95227,
  75.41367,
  -53.64331,
  75.37709,
  -54.16016,
  75.40265,
  -54.49108,
  75.405,
  -53.29064,
  75.43598,
  -53.27973,
  75.55351,
  -53.97705,
  75.35275,
  -54.53227,
  75.26194,
  -54.41441,
  75.51382,
  -53.25823,
  75.53917,
  -53.67912,
  75.32951,
  -54.31174,
  75.39924,
  -54.6587,
  75.35934,
  -53.83406,
  75.42509,
  -53.57505,
  75.42735,
  -54.31968,
  75.50877,
  -54.77357,
  75.3229,
  -54.737,
  75.36761,
  -53.98958,
  75.47401,
  -53.83375,
  75.48244,
  -54.4837,
  75.22174,
  -54.77822,
  75.22047,
  -54.5752,
  75.49251,
  -53.80748,
  75.44043,
  -54.33756,
  75.3713,
  -54.68293,
  75.08734,
  -54.84767,
  75.24926,
  -54.74097,
  75.44522,
  -54.16355,
  75.34815,
  -54.69554,
  75.20778,
  -55.18597,
  75.26942,
  -55.25907,
  75.41686,
  -53.98673,
  75.40319,
  -54.46646,
  75.33168,
  -54.97514,
  75.22417,
  -55.08517,
  75.30054,
  -53.92952,
  75.52354,
  -54.14849,
  75.46046,
  -54.74057,
  75.25597,
  -55.12278,
  75.2781,
  -53.70147,
  75.4632,
  -53.84176,
  75.36569,
  -54.47032,
  75.2555,
  -54.80178,
  75.48221,
  -53.31939,
  75.5262,
  -53.7253,
  75.52844,
  -54.26201,
  75.19355,
  -54.77756,
  75.31026,
  -53.63806,
  75.36691,
  -53.46946,
  75.58596,
  -54.0078,
  75.29647,
  -54.51898,
  75.21104,
  -54.4077,
  75.48537,
  -53.46729,
  75.5023,
  -53.93951,
  75.20886,
  -54.46327,
  75.17556,
  -54.51845,
  75.37657,
  -54.26071,
  75.47525,
  -53.72545,
  75.39117,
  -54.21247,
  75.39406,
  -54.56694,
  75.30214,
  -54.39057,
  75.18605,
  -53.80988,
  75.24158,
  -54.45673,
  75.28667,
  -54.56109,
  75.21368,
  -54.58276,
  75.33286,
  -54.18266,
  75.40226,
  -54.24049,
  75.3411,
  -54.38681,
  75.25465,
  -54.84959,
  75.22734,
  -54.39397,
  75.41729,
  -54.11338,
  75.43217,
  -54.14319,
  75.33526,
  -54.74945,
  75.18126,
  -55.28876,
  75.25134,
  -54.3506,
  75.33007,
  -54.06221,
  75.38367,
  -54.58786,
  75.22655,
  -55.14116,
  75.26866,
  -55.26443,
  75.30442,
  -54.03084,
  75.50806,
  -54.10094,
  75.31098,
  -54.76185,
  75.16203,
  -55.2462,
  75.34579,
  -53.96214,
  75.44284,
  -54.07473,
  75.23129,
  -54.55927,
  75.16217,
  -54.91403,
  75.24778,
  -53.61563,
  75.38491,
  -53.64509,
  75.37368,
  -54.47743,
  75.45118,
  -54.93583,
  75.39223,
  -54.15773,
  75.44263,
  -53.53554,
  75.28578,
  -54.05236,
  75.4323,
  -54.61211,
  75.42654,
  -53.9291,
  75.43514,
  -53.67169,
  75.35548,
  -54.11614,
  75.31292,
  -54.33876,
  75.3387,
  -54.20326,
  75.29365,
  -53.43858,
  75.39999,
  -53.57924,
  75.36909,
  -54.14893,
  75.17276,
  -54.76834,
  75.34224,
  -53.64019,
  75.50484,
  -53.60596,
  75.24625,
  -54.56942,
  75.22095,
  -54.61148,
  75.29385,
  -54.72705,
  75.19127,
  -53.99551,
  75.44002,
  -53.89434,
  75.44141,
  -54.35485,
  75.31389,
  -54.74089,
  75.25904,
  -54.57575,
  75.29982,
  -54.36477,
  75.38258,
  -54.33023,
  75.30313,
  -54.6627,
  75.30887,
  -55.04218,
  75.32429,
  -54.72547,
  75.35476,
  -54.17981,
  75.45914,
  -54.28037,
  75.26644,
  -54.76948,
  75.32586,
  -54.67377,
  75.32284,
  -54.19804,
  75.55959,
  -54.1589,
  75.37524,
  -54.78408,
  75.14333,
  -55.13877,
  75.43851,
  -54.02288,
  75.42819,
  -53.97285,
  75.37698,
  -54.48059,
  75.22236,
  -55.08588,
  75.17551,
  -54.0709,
  75.4743,
  -53.68643,
  75.38226,
  -54.37297,
  75.28922,
  -54.82468,
  75.25927,
  -53.79391,
  75.55649,
  -53.5075,
  75.41096,
  -54.07007,
  75.29647,
  -54.62543,
  75.42217,
  -53.9098,
  75.396,
  -53.40115,
  75.4903,
  -53.859,
  75.4784,
  -54.4495,
  75.27647,
  -54.44284,
  75.33399,
  -53.40657,
  75.42719,
  -53.66221,
  -14.22611,
  -77.68449,
  -14.66727,
  -77.65236,
  -13.57793,
  -77.18984,
  -13.94214,
  -77.56248,
  -14.28421,
  -77.55075,
  -14.55616,
  -77.62982,
  -13.86991,
  -77.3364,
  -14.3271,
  -77.6385,
  -14.1154,
  -77.65112,
  -14.71269,
  -77.76078,
  -14.50649,
  -77.6638,
  -15.17249,
  -77.89623,
  -14.32831,
  -77.50005,
  -14.4868,
  -77.81565,
  -15.17351,
  -77.88645,
  -14.14832,
  -77.3691,
  -13.79397,
  -77.50333,
  -14.49368,
  -77.65751,
  -14.60266,
  -77.56497,
  -14.22078,
  -77.4825,
  -14.13271,
  -77.4537,
  -14.19472,
  -77.50739,
  -13.48724,
  -77.26214,
  -13.9379,
  -77.49413,
  -14.61808,
  -77.79191,
  -14.32246,
  -77.56191,
  -14.49095,
  -77.58853,
  -14.36612,
  -77.58026,
  -15.19823,
  -77.77856,
  -14.2,
  -77.51107,
  -14.62934,
  -77.712,
  -15.2589,
  -77.90833,
  -14.69009,
  -77.63795,
  -13.94278,
  -77.59393,
  -14.48192,
  -77.76381,
  -14.64612,
  -77.52103,
  -13.46911,
  -77.20545,
  -14.03464,
  -77.48817,
  -14.25383,
  -77.70805,
  -13.82867,
  -77.36057,
  -13.73678,
  -77.40066,
  -13.68545,
  -77.42338,
  -14.20706,
  -77.59487,
  -14.71686,
  -77.68497,
  -15.03693,
  -77.81213,
  -14.88661,
  -77.71411,
  -14.27692,
  -77.53953,
  -14.50965,
  -77.7781,
  -15.20689,
  -77.85256,
  -15.36814,
  -77.85546,
  -14.05969,
  -77.3513,
  -14.45578,
  -77.6188,
  -14.98228,
  -77.86124,
  -14.94745,
  -77.72793,
  -13.68428,
  -77.42947,
  -14.15347,
  -77.69764,
  -14.79527,
  -77.68385,
  -13.89116,
  -77.29482,
  -14.10654,
  -77.5601,
  -14.09988,
  -77.52631,
  -14.22511,
  -77.61697,
  -14.33797,
  -77.69594,
  -14.71953,
  -77.63065,
  -14.16238,
  -77.39089,
  -14.30371,
  -77.75222,
  -14.65292,
  -77.67383,
  -14.97735,
  -77.82304,
  -14.85907,
  -77.86018,
  -14.52167,
  -77.61987,
  -14.76522,
  -77.79738,
  -15.35681,
  -77.97124,
  -14.94682,
  -77.64253,
  -13.9871,
  -77.60714,
  -14.62699,
  -77.7142,
  -15.19583,
  -77.9387,
  -14.1533,
  -77.34686,
  -13.88076,
  -77.42064,
  -14.46014,
  -77.60462,
  -14.87263,
  -77.77522,
  -14.03466,
  -77.41019,
  -13.83355,
  -77.31379,
  -14.2051,
  -77.65916,
  -14.67204,
  -77.87844,
  -14.529,
  -77.55229,
  -13.78591,
  -77.29118,
  -13.90053,
  -77.56076,
  -14.06005,
  -77.52517,
  -14.85007,
  -77.77479,
  -14.98165,
  -77.68703,
  -14.15705,
  -77.4623,
  -14.35436,
  -77.60439,
  -14.68948,
  -77.7961,
  -15.33887,
  -77.95439,
  -14.74068,
  -77.68169,
  -14.34758,
  -77.67397,
  -14.88284,
  -77.8671,
  -15.39357,
  -78.03759,
  -14.77388,
  -77.63039,
  -14.06666,
  -77.41568,
  -14.55172,
  -77.74725,
  -15.18549,
  -77.8911,
  -14.72207,
  -77.53986,
  -13.88165,
  -77.46487,
  -14.35905,
  -77.72398,
  -14.98699,
  -77.80529,
  -14.03429,
  -77.37096,
  -13.6721,
  -77.33815,
  -14.23597,
  -77.59033,
  -14.70746,
  -77.81149,
  -14.63099,
  -77.71947,
  -13.76768,
  -77.33231,
  -14.0347,
  -77.5126,
  -14.47381,
  -77.71764,
  -14.72417,
  -77.72462,
  -14.50563,
  -77.55444,
  -13.8311,
  -77.45905,
  -14.2625,
  -77.67675,
  -14.89499,
  -77.74629,
  -15.30678,
  -77.8987,
  -14.57711,
  -77.58272,
  -14.12513,
  -77.57543,
  -14.47426,
  -77.56287,
  -15.27161,
  -77.95246,
  -15.57284,
  -77.92033,
  -14.71881,
  -77.59734,
  -14.54914,
  -77.74187,
  -14.91743,
  -77.84224,
  -15.13446,
  -77.93935,
  -14.18128,
  -77.34209,
  -14.29475,
  -77.65765,
  -14.76143,
  -77.8592,
  -15.39743,
  -77.81184,
  -14.17025,
  -77.28748,
  -13.96128,
  -77.50477,
  -14.63412,
  -77.68224,
  -15.16452,
  -77.76639,
  -14.32976,
  -77.42674,
  -13.90117,
  -77.40836,
  -14.42609,
  -77.55147,
  -14.97586,
  -77.78011,
  -14.16573,
  -77.35449,
  -13.83263,
  -77.34474,
  -14.15437,
  -77.56757,
  -14.67096,
  -77.66588,
  -13.72817,
  -77.2532,
  -13.52717,
  -77.27648,
  -14.05219,
  -77.62422,
  -14.45814,
  -77.7288,
  -14.99055,
  -77.82172,
  -14.38631,
  -77.51278,
  -13.89222,
  -77.52826,
  -14.48354,
  -77.72324,
  -14.6524,
  -77.7233,
  -14.88101,
  -77.78097,
  -14.3807,
  -77.58812,
  -14.02726,
  -77.54978,
  -14.64667,
  -77.83348,
  -15.29493,
  -77.97856,
  -15.64287,
  -77.92805,
  -14.54764,
  -77.61349,
  -14.56869,
  -77.71014,
  -14.97384,
  -77.92414,
  -15.43881,
  -77.96307,
  -14.48502,
  -77.47847,
  -14.21796,
  -77.71436,
  -14.73209,
  -77.79946,
  -15.2102,
  -77.9033,
  -14.23137,
  -77.52467,
  -13.80445,
  -77.62361,
  -14.64684,
  -77.71798,
  -15.16628,
  -77.83173,
  -14.16367,
  -77.36317,
  -13.85869,
  -77.29453,
  -14.36021,
  -77.61031,
  -14.71011,
  -77.79643,
  -13.58733,
  -77.2123,
  -13.65087,
  -77.25578,
  -14.11759,
  -77.61141,
  -14.64799,
  -77.82405,
  -14.622,
  -77.59319,
  -13.50153,
  -77.2692,
  -13.92234,
  -77.46346,
  -14.50523,
  -77.64779,
  -14.79593,
  -77.80107,
  -14.06598,
  -77.4876,
  -13.87332,
  -77.30879,
  -14.51872,
  -77.74992,
  -14.85273,
  -77.82487,
  -14.85309,
  -77.7072,
  -14.29099,
  -77.51287,
  -14.07456,
  -77.54951,
  -14.57912,
  -77.77957,
  -14.96981,
  -77.73344,
  -14.83262,
  -77.56297,
  -14.06875,
  -77.49812,
  -14.50031,
  -77.6908,
  -14.79816,
  -77.83287,
  -15.01328,
  -77.65139,
  -14.93933,
  -77.67889,
  -14.29445,
  -77.62045,
  -14.86765,
  -77.74445,
  -15.31992,
  -77.95836,
  -15.39163,
  -78.01579,
  -14.15027,
  -77.52728,
  -14.59214,
  -77.74561,
  -15.10115,
  -77.94356,
  -15.29973,
  -77.87025,
  -14.16257,
  -77.36768,
  -14.26119,
  -77.71517,
  -14.85956,
  -77.93626,
  -15.26915,
  -77.76627,
  -13.97507,
  -77.28825,
  -14.02236,
  -77.61825,
  -14.66078,
  -77.70556,
  -14.9743,
  -77.74224,
  -13.45524,
  -77.28119,
  -13.93555,
  -77.56461,
  -14.50039,
  -77.65386,
  -14.95632,
  -77.80871,
  -13.93687,
  -77.32011,
  -13.80009,
  -77.21938,
  -14.18596,
  -77.72627,
  -14.68249,
  -77.78151,
  -14.6285,
  -77.60478,
  -13.71599,
  -77.29681,
  -14.06586,
  -77.55463,
  -14.62166,
  -77.66806,
  -14.74049,
  -77.78249,
  -14.4505,
  -77.59968,
  -13.93995,
  -77.41051,
  -14.33845,
  -77.60042,
  -14.80618,
  -77.75087,
  -14.65256,
  -77.62537,
  -14.11147,
  -77.25368,
  -14.48204,
  -77.64352,
  -14.71348,
  -77.6834,
  -14.81606,
  -77.6571,
  -14.46154,
  -77.58753,
  -14.42583,
  -77.55718,
  -14.67533,
  -77.58926,
  -15.00728,
  -77.7762,
  -14.58295,
  -77.68156,
  -14.32835,
  -77.58721,
  -14.28408,
  -77.65067,
  -14.89589,
  -77.79637,
  -15.31974,
  -77.90044,
  -14.47767,
  -77.5695,
  -14.22492,
  -77.48806,
  -14.74257,
  -77.61623,
  -15.30886,
  -78.04389,
  -15.23856,
  -77.95309,
  -14.14418,
  -77.48399,
  -14.26879,
  -77.66641,
  -15.11452,
  -77.74654,
  -15.46572,
  -77.95094,
  -14.18366,
  -77.45116,
  -14.20384,
  -77.67905,
  -14.82109,
  -77.66947,
  -15.12344,
  -77.76174,
  -13.94865,
  -77.20683,
  -13.93399,
  -77.41659,
  -14.55163,
  -77.75021,
  -14.96032,
  -77.96703,
  -14.32241,
  -77.55685,
  -13.81945,
  -77.32147,
  -14.33341,
  -77.57384,
  -14.70792,
  -77.71756,
  -14.35042,
  -77.52592,
  -13.83475,
  -77.29808,
  -14.32437,
  -77.54939,
  -14.55144,
  -77.60152,
  -14.44692,
  -77.53131,
  -13.6795,
  -77.15056,
  -13.8709,
  -77.41315,
  -14.29999,
  -77.67805,
  -14.91482,
  -77.78239,
  -13.85426,
  -77.31986,
  -13.80914,
  -77.38786,
  -14.77996,
  -77.66796,
  -14.80933,
  -77.6172,
  -14.92895,
  -77.78773,
  -14.31943,
  -77.33208,
  -14.05001,
  -77.44673,
  -14.53109,
  -77.75127,
  -14.89514,
  -77.86423,
  -14.77049,
  -77.71277,
  -14.60507,
  -77.62816,
  -14.50844,
  -77.65356,
  -14.8162,
  -77.79929,
  -15.16681,
  -77.96514,
  -14.86382,
  -77.75005,
  -14.30791,
  -77.54717,
  -14.44137,
  -77.74139,
  -14.88562,
  -77.82546,
  -14.82699,
  -77.80572,
  -14.35464,
  -77.42073,
  -14.16449,
  -77.68037,
  -14.85523,
  -77.87627,
  -15.28118,
  -77.91873,
  -14.1748,
  -77.55824,
  -14.13898,
  -77.56207,
  -14.68475,
  -77.75585,
  -15.26102,
  -77.82855,
  -14.34724,
  -77.35941,
  -13.91392,
  -77.42021,
  -14.44816,
  -77.67558,
  -14.95393,
  -77.77574,
  -14.07017,
  -77.24312,
  -13.68025,
  -77.39658,
  -14.23736,
  -77.60903,
  -14.87104,
  -77.78573,
  -14.11498,
  -77.42229,
  -13.64874,
  -77.22375,
  -14.03749,
  -77.54807,
  -14.53753,
  -77.74079,
  -14.62295,
  -77.64018,
  -13.69655,
  -77.15564,
  -13.89584,
  -77.37731,
  -65.4136,
  -17.31545,
  -65.66879,
  -16.86457,
  -64.67429,
  -17.64606,
  -65.14156,
  -17.5406,
  -65.36923,
  -17.17989,
  -65.61687,
  -17.00402,
  -65.02346,
  -17.5443,
  -65.43049,
  -17.22604,
  -65.31678,
  -17.40587,
  -65.79259,
  -16.89435,
  -65.51939,
  -16.99392,
  -65.98582,
  -16.56401,
  -65.34724,
  -17.16081,
  -65.67336,
  -17.17053,
  -66.09493,
  -16.52214,
  -65.15239,
  -17.22781,
  -65.13319,
  -17.62809,
  -65.6367,
  -17.1291,
  -65.59461,
  -16.98622,
  -65.24038,
  -17.12525,
  -65.07199,
  -17.30094,
  -65.36268,
  -17.26891,
  -64.68094,
  -17.76766,
  -65.16306,
  -17.4185,
  -65.70817,
  -17.05151,
  -65.54395,
  -17.2228,
  -65.47012,
  -17.04599,
  -65.41509,
  -17.21678,
  -66.05148,
  -16.53701,
  -65.28555,
  -17.37264,
  -65.72754,
  -17.06043,
  -66.15897,
  -16.55838,
  -65.54787,
  -16.95716,
  -65.16622,
  -17.54364,
  -65.59259,
  -17.11258,
  -65.53957,
  -16.87813,
  -64.5818,
  -17.73322,
  -65.1082,
  -17.45738,
  -65.42698,
  -17.35717,
  -64.91531,
  -17.51686,
  -64.94831,
  -17.64612,
  -64.97105,
  -17.69325,
  -65.29108,
  -17.33554,
  -65.73941,
  -16.9185,
  -66.02723,
  -16.57476,
  -65.69793,
  -16.80672,
  -65.35004,
  -17.24775,
  -65.71232,
  -17.19592,
  -66.14458,
  -16.64243,
  -66.08742,
  -16.45742,
  -65.05412,
  -17.3876,
  -65.50035,
  -17.14974,
  -65.8932,
  -16.8185,
  -65.66531,
  -16.77991,
  -64.91454,
  -17.70176,
  -65.36417,
  -17.4383,
  -65.65968,
  -16.928,
  -64.92522,
  -17.45603,
  -65.16066,
  -17.36914,
  -65.17289,
  -17.37957,
  -65.29445,
  -17.31087,
  -65.42591,
  -17.24259,
  -65.59834,
  -16.90846,
  -65.0518,
  -17.31906,
  -65.56509,
  -17.27248,
  -65.61161,
  -17.02073,
  -65.80602,
  -16.7756,
  -65.84576,
  -16.85386,
  -65.48976,
  -17.15793,
  -65.77794,
  -16.94801,
  -66.22222,
  -16.54594,
  -65.69975,
  -16.7118,
  -65.19217,
  -17.52367,
  -65.71246,
  -16.99064,
  -66.14365,
  -16.56097,
  -65.0961,
  -17.25074,
  -65.07049,
  -17.52748,
  -65.53711,
  -17.12208,
  -65.84769,
  -16.78749,
  -65.13745,
  -17.24428,
  -64.8541,
  -17.46768,
  -65.49252,
  -17.34868,
  -65.80704,
  -17.07225,
  -65.47779,
  -17.06184,
  -64.90906,
  -17.62169,
  -65.36239,
  -17.52216,
  -65.23944,
  -17.36934,
  -65.87533,
  -16.86575,
  -65.79723,
  -16.68737,
  -65.25683,
  -17.29705,
  -65.45023,
  -17.19605,
  -65.73119,
  -17.16815,
  -66.20834,
  -16.48936,
  -65.63289,
  -16.90127,
  -65.43767,
  -17.21124,
  -65.80921,
  -16.85065,
  -66.26577,
  -16.50797,
  -65.65154,
  -16.7652,
  -65.15229,
  -17.35793,
  -65.58071,
  -17.05051,
  -66.06771,
  -16.62245,
  -65.4465,
  -16.88117,
  -64.9891,
  -17.56809,
  -65.56495,
  -17.24459,
  -65.89011,
  -16.73516,
  -65.03742,
  -17.44224,
  -64.84667,
  -17.79194,
  -65.36618,
  -17.33582,
  -65.87181,
  -16.91163,
  -65.6152,
  -17.01048,
  -64.80544,
  -17.53041,
  -65.11933,
  -17.39159,
  -65.54987,
  -17.14266,
  -65.67567,
  -16.93864,
  -65.4463,
  -16.9363,
  -65.06026,
  -17.50682,
  -65.5189,
  -17.29402,
  -65.80636,
  -16.91574,
  -66.06483,
  -16.49912,
  -65.53575,
  -16.92817,
  -65.28113,
  -17.32918,
  -65.53261,
  -17.1174,
  -66.21879,
  -16.63403,
  -66.34425,
  -16.27964,
  -65.66501,
  -16.93845,
  -65.56926,
  -16.97583,
  -65.939,
  -16.7079,
  -66.02677,
  -16.57191,
  -65.04559,
  -17.21778,
  -65.2891,
  -17.36287,
  -65.80398,
  -16.94683,
  -66.14074,
  -16.37448,
  -65.06702,
  -17.1872,
  -65.23199,
  -17.50333,
  -65.60998,
  -16.99762,
  -65.93317,
  -16.53249,
  -65.19358,
  -17.09374,
  -64.98878,
  -17.56582,
  -65.48833,
  -17.18112,
  -65.8596,
  -16.7384,
  -65.14354,
  -17.21918,
  -64.92284,
  -17.56188,
  -65.30698,
  -17.29184,
  -65.71272,
  -16.96788,
  -64.85424,
  -17.57573,
  -64.69997,
  -17.73363,
  -65.25862,
  -17.49399,
  -65.59097,
  -17.1166,
  -65.8697,
  -16.82237,
  -65.3186,
  -17.10605,
  -65.13284,
  -17.50175,
  -65.52362,
  -17.20177,
  -65.71736,
  -17.0102,
  -65.81969,
  -16.768,
  -65.38956,
  -17.11209,
  -65.3202,
  -17.45334,
  -65.73111,
  -17.02074,
  -66.14649,
  -16.61606,
  -66.36336,
  -16.35251,
  -65.61518,
  -17.09956,
  -65.63387,
  -17.04305,
  -65.99941,
  -16.87428,
  -66.25779,
  -16.43367,
  -65.32607,
  -16.94483,
  -65.28927,
  -17.28366,
  -65.8113,
  -16.87819,
  -66.07552,
  -16.55594,
  -65.25752,
  -17.32905,
  -65.21776,
  -17.55762,
  -65.68289,
  -17.02563,
  -66.0263,
  -16.67901,
  -65.24593,
  -17.24352,
  -64.99786,
  -17.53933,
  -65.55932,
  -17.20984,
  -65.70011,
  -17.02349,
  -64.72225,
  -17.67297,
  -64.65107,
  -17.69513,
  -65.34717,
  -17.4549,
  -65.70824,
  -17.01204,
  -65.48903,
  -17.00043,
  -64.70119,
  -17.77437,
  -65.11494,
  -17.56878,
  -65.57893,
  -17.06824,
  -65.84303,
  -16.93047,
  -65.15114,
  -17.43583,
  -64.90158,
  -17.55132,
  -65.60751,
  -17.19142,
  -65.93345,
  -16.90702,
  -65.7959,
  -16.84223,
  -65.30917,
  -17.23953,
  -65.19015,
  -17.39762,
  -65.68808,
  -17.07271,
  -65.89011,
  -16.7203,
  -65.73384,
  -16.78081,
  -65.18789,
  -17.4627,
  -65.48322,
  -17.17061,
  -65.89466,
  -16.91747,
  -65.82989,
  -16.70115,
  -65.79685,
  -16.6877,
  -65.43296,
  -17.19184,
  -65.79544,
  -16.84646,
  -66.20834,
  -16.44394,
  -66.25231,
  -16.47211,
  -65.31441,
  -17.30787,
  -65.64532,
  -17.07093,
  -66.04717,
  -16.75897,
  -66.11391,
  -16.5124,
  -65.09577,
  -17.27048,
  -65.42595,
  -17.33057,
  -65.92611,
  -16.88039,
  -66.1107,
  -16.53036,
  -64.94862,
  -17.42986,
  -65.32838,
  -17.54066,
  -65.69572,
  -17.01096,
  -65.92395,
  -16.61395,
  -64.67792,
  -17.71678,
  -65.12124,
  -17.52883,
  -65.52708,
  -17.25541,
  -65.86211,
  -16.82232,
  -64.96172,
  -17.38801,
  -64.81756,
  -17.59214,
  -65.3383,
  -17.36878,
  -65.70287,
  -17.07122,
  -65.52787,
  -16.93734,
  -64.84846,
  -17.66766,
  -65.2864,
  -17.42506,
  -65.63422,
  -17.03601,
  -65.71009,
  -16.79371,
  -65.4334,
  -17.09656,
  -65.0999,
  -17.38993,
  -65.55564,
  -17.21666,
  -65.81474,
  -16.94444,
  -65.5048,
  -17.01373,
  -65.00552,
  -17.33883,
  -65.6601,
  -16.93491,
  -65.66124,
  -16.7982,
  -65.65498,
  -16.75309,
  -65.43763,
  -17.0482,
  -65.52513,
  -17.10456,
  -65.60825,
  -16.98089,
  -65.88806,
  -16.70184,
  -65.47815,
  -16.92927,
  -65.40737,
  -17.12625,
  -65.42101,
  -17.22795,
  -65.81525,
  -16.82844,
  -66.15499,
  -16.46707,
  -65.66698,
  -17.02043,
  -65.22378,
  -17.2444,
  -65.71648,
  -16.90278,
  -66.21609,
  -16.59329,
  -66.2047,
  -16.51548,
  -65.17854,
  -17.28729,
  -65.50632,
  -17.3997,
  -65.96799,
  -16.90122,
  -66.2174,
  -16.42444,
  -65.1788,
  -17.24247,
  -65.43721,
  -17.34045,
  -65.69265,
  -16.82738,
  -65.96646,
  -16.59011,
  -64.84525,
  -17.28774,
  -65.06837,
  -17.49044,
  -65.63849,
  -17.08027,
  -66.04486,
  -16.82393,
  -65.3046,
  -17.20261,
  -64.91376,
  -17.57021,
  -65.43085,
  -17.27434,
  -65.74316,
  -16.83323,
  -65.22941,
  -17.25269,
  -64.91863,
  -17.53299,
  -65.27059,
  -17.20961,
  -65.53589,
  -17.02228,
  -65.45172,
  -17.14399,
  -64.70564,
  -17.53323,
  -64.93234,
  -17.52777,
  -65.40356,
  -17.27291,
  -65.7463,
  -16.81972,
  -64.94446,
  -17.54501,
  -64.9896,
  -17.57903,
  -65.65927,
  -16.86263,
  -65.66424,
  -16.79192,
  -65.85395,
  -16.86788,
  -65.11132,
  -17.14472,
  -65.13326,
  -17.43316,
  -65.6098,
  -17.18105,
  -65.99287,
  -16.81831,
  -65.69089,
  -16.87596,
  -65.55578,
  -17.01327,
  -65.51942,
  -17.11365,
  -65.77191,
  -16.84866,
  -66.03346,
  -16.62074,
  -65.81143,
  -16.80344,
  -65.39483,
  -17.2298,
  -65.56667,
  -17.11049,
  -65.87546,
  -16.78226,
  -65.81636,
  -16.86609,
  -65.26316,
  -17.15839,
  -65.43443,
  -17.31758,
  -65.85508,
  -16.88068,
  -66.06793,
  -16.57218,
  -65.21304,
  -17.31335,
  -65.21503,
  -17.34257,
  -65.70286,
  -17.01162,
  -66.12071,
  -16.57997,
  -65.1683,
  -17.06827,
  -65.10743,
  -17.47272,
  -65.5929,
  -17.11454,
  -65.86874,
  -16.78018,
  -64.96012,
  -17.31385,
  -64.92161,
  -17.65481,
  -65.3351,
  -17.1768,
  -65.81267,
  -16.82844,
  -65.19736,
  -17.30173,
  -64.74113,
  -17.70844,
  -65.2647,
  -17.44154,
  -65.65023,
  -17.07519,
  -65.54909,
  -17.01077,
  -64.68964,
  -17.55024,
  -65.0283,
  -17.5191 ;

 jsrc_mask =
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1,
  1 ;

 sigma_c = 4.567846, 4.568751, 4.5683, 4.569418, 4.56914, 4.57147, 4.579232, 
    4.579414, 4.575336, 4.574708, 4.573055, 4.57149, 4.573745, 4.576893, 
    4.58806, 4.592668, 4.581561, 4.570082, 4.564, 4.561146, 4.564439, 
    4.562511, 4.557363, 4.5597, 4.563426, 4.566694, 4.5675, 4.568791, 
    4.569862, 4.571967, 4.571446, 4.573476, 4.573061, 4.570632, 4.568616, 
    4.578717, 4.593209, 4.612979, 4.618958, 4.621602, 4.630395, 4.639049, 
    4.6397, 4.6394, 4.630472, 4.622649, 4.617032, 4.61768, 4.609563, 
    4.594225, 4.597661, 4.602603, 4.616725, 4.623173, 4.612912, 4.611436, 
    4.631897, 4.634503, 4.6336, 4.624523, 4.595595, 4.588931, 4.588986, 
    4.587251, 4.588737, 4.596098, 4.621344, 4.629237, 4.624228, 4.61436, 
    4.615736, 4.617553, 4.617139, 4.624625, 4.6251, 4.625546, 4.613909, 
    4.60956, 4.614627, 4.607135, 4.612123, 4.59813, 4.600029, 4.611267, 
    4.602, 4.60034, 4.605921, 4.604317, 4.608295, 4.607721, 4.606894, 
    4.608646, 4.611225, 4.614689, 4.610782, 4.610355, 4.610455, 4.611791, 
    4.611824, 4.612126, 4.61374, 4.614515, 4.600904, 4.616194, 4.617256, 
    4.618858, 4.617721, 4.6166, 4.616983, 4.617316, 4.617379, 4.6173, 4.6175, 
    4.617187, 4.617701, 4.618, 4.617566, 4.616617, 4.617313, 4.61707, 4.6173, 
    4.61785, 4.6179, 4.618523, 4.619482, 4.6201, 4.619843, 4.618685, 
    4.620242, 4.622736, 4.622365, 4.6218, 4.622515, 4.627153, 4.624638, 
    4.629638, 4.633592, 4.634627, 4.621542, 4.62545, 4.623494, 4.621653, 
    4.626216, 4.633325, 4.632357, 4.63609, 4.639235, 4.62957, 4.626738, 
    4.630363, 4.631992, 4.621841, 4.624331, 4.627941, 4.626648, 4.626985, 
    4.624753, 4.624873, 4.625373, 4.62459, 4.622435, 4.622191, 4.623002, 
    4.624955, 4.627852, 4.625674, 4.620615, 4.620259, 4.617554, 4.619176, 
    4.623729, 4.617635, 4.628175, 4.618324, 4.619489, 4.6216, 4.621587, 
    4.622174, 4.622208, 4.622389, 4.624587, 4.626148, 4.62562, 4.623461, 
    4.623142, 4.622468, 4.622107, 4.622366, 4.621219, 4.622059, 4.621865, 
    4.62261, 4.622975, 4.62321, 4.622665, 4.622643, 4.622592, 4.622547, 
    4.62307, 4.623375, 4.621956, 4.621641, 4.6193, 4.622584, 4.623941, 
    4.624394, 4.6249, 4.624731, 4.637477, 4.625443, 4.625505, 4.623164, 
    4.621059, 4.61907, 4.622075, 4.642486, 4.647761, 4.648807, 4.64808, 
    4.636666, 4.621532, 4.610478, 4.621891, 4.631329, 4.646948, 4.647325, 
    4.614202, 4.609656, 4.61023, 4.610591, 4.609763, 4.6109, 4.632373, 
    4.641195, 4.64444, 4.641116, 4.622263, 4.611711, 4.611494, 4.612621, 
    4.613647, 4.614656, 4.641466, 4.64132, 4.638702, 4.634595, 4.618063, 
    4.594851, 4.576742, 4.582653, 4.610582, 4.619941, 4.622076, 4.624018, 
    4.624214, 4.622211, 4.621377, 4.609036, 4.586376, 4.582213, 4.585155, 
    4.59831, 4.615165, 4.607287, 4.611683, 4.600698, 4.601643, 4.629858, 
    4.630089, 4.634055, 4.633235, 4.629064, 4.629391, 4.624741, 4.604583, 
    4.620414, 4.628816, 4.620861, 4.627119, 4.632283, 4.62801, 4.618903, 
    4.627518, 4.633946, 4.63526, 4.642232, 4.642746, 4.643812, 4.642117, 
    4.638324, 4.637309, 4.635895, 4.634771, 4.617516, 4.627507, 4.62509, 
    4.638824, 4.636388, 4.627536, 4.639615, 4.646664, 4.629085, 4.609486, 
    4.609216, 4.614288, 4.63878, 4.623609, 4.61618, 4.617441, 4.639076, 
    4.637013, 4.642406, 4.661279, 4.665342, 4.657032, 4.625436, 4.629019, 
    4.6355 ;

 time =
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26,
  1295253367.44, 1295253528.68,
  1295253367.44, 1295253528.68,
  1295253444.96, 1295253606.2,
  1295253444.96, 1295253606.2,
  1295253523.12, 1295253684.36,
  1295253523.12, 1295253684.36,
  1295253600.34, 1295253761.58,
  1295253600.34, 1295253761.58,
  1295253678.4, 1295253839.64,
  1295253678.4, 1295253839.64,
  1295253756.08, 1295253917.32,
  1295253756.08, 1295253917.32,
  1295253832.84, 1295253994.08,
  1295253832.84, 1295253994.08,
  1295253910.96, 1295254072.2,
  1295253910.96, 1295254072.2,
  1295253988.86, 1295254150.1,
  1295253988.86, 1295254150.1,
  1295254067.02, 1295254228.26,
  1295254067.02, 1295254228.26,
  1295254145.28, 1295254306.52,
  1295254145.28, 1295254306.52,
  1295254222.7, 1295254383.94,
  1295254222.7, 1295254383.94,
  1295254299.8, 1295254461.04,
  1295254299.8, 1295254461.04,
  1295254377.5, 1295254538.74,
  1295254377.5, 1295254538.74,
  1295254454.8, 1295254616.04,
  1295254454.8, 1295254616.04,
  1295254532.74, 1295254693.98,
  1295254532.74, 1295254693.98,
  1295254611.42, 1295254772.66,
  1295254611.42, 1295254772.66,
  1295254689.66, 1295254850.9,
  1295254689.66, 1295254850.9,
  1295254767.84, 1295254929.08,
  1295254767.84, 1295254929.08,
  1295254844.68, 1295255005.92,
  1295254844.68, 1295255005.92,
  1295254923.06, 1295255084.3,
  1295254923.06, 1295255084.3,
  1295255001.22, 1295255162.46,
  1295255001.22, 1295255162.46,
  1295255078.68, 1295255239.92,
  1295255078.68, 1295255239.92,
  1295255156.32, 1295255317.56,
  1295255156.32, 1295255317.56,
  1295255233.96, 1295255395.2,
  1295255233.96, 1295255395.2,
  1295255311.76, 1295255473,
  1295255311.76, 1295255473,
  1295255389.6, 1295255550.84,
  1295255389.6, 1295255550.84,
  1295255467.16, 1295255628.4,
  1295255467.16, 1295255628.4,
  1295255544.36, 1295255705.6,
  1295255544.36, 1295255705.6,
  1295255622.62, 1295255783.86,
  1295255622.62, 1295255783.86,
  1295255700.86, 1295255862.1,
  1295255700.86, 1295255862.1,
  1295255779.28, 1295255940.52,
  1295255779.28, 1295255940.52,
  1295255856.4, 1295256017.64,
  1295255856.4, 1295256017.64,
  1295255934.64, 1295256095.88,
  1295255934.64, 1295256095.88,
  1295256011.58, 1295256172.82,
  1295256011.58, 1295256172.82,
  1295256089.6, 1295256250.84,
  1295256089.6, 1295256250.84,
  1295256166.32, 1295256327.56,
  1295256166.32, 1295256327.56,
  1295256243.76, 1295256405,
  1295256243.76, 1295256405,
  1295256321.86, 1295256483.1,
  1295256321.86, 1295256483.1,
  1295256399.1, 1295256560.34,
  1295256399.1, 1295256560.34,
  1295256477.14, 1295256638.38,
  1295256477.14, 1295256638.38,
  1295256554.8, 1295256716.04,
  1295256554.8, 1295256716.04,
  1295256632.46, 1295256793.7,
  1295256632.46, 1295256793.7,
  1295256710.16, 1295256871.4,
  1295256710.16, 1295256871.4,
  1295256788.14, 1295256949.38,
  1295256788.14, 1295256949.38,
  1295256866.28, 1295257027.52,
  1295256866.28, 1295257027.52,
  1295256943.58, 1295257104.82,
  1295256943.58, 1295257104.82,
  1295257020.38, 1295257181.62,
  1295257020.38, 1295257181.62,
  1295257098.28, 1295257259.52,
  1295257098.28, 1295257259.52,
  1295257176.06, 1295257337.3,
  1295257176.06, 1295257337.3,
  1295257254.08, 1295257415.32,
  1295257254.08, 1295257415.32,
  1295257332.24, 1295257493.48,
  1295257332.24, 1295257493.48,
  1295257410.52, 1295257571.76,
  1295257410.52, 1295257571.76,
  1295257488.44, 1295257649.68,
  1295257488.44, 1295257649.68,
  1295257566.96, 1295257728.2,
  1295257566.96, 1295257728.2,
  1295257645.1, 1295257806.34,
  1295257645.1, 1295257806.34,
  1295257722.42, 1295257883.66,
  1295257722.42, 1295257883.66,
  1295257800.76, 1295257962,
  1295257800.76, 1295257962,
  1295257879, 1295258040.24,
  1295257879, 1295258040.24,
  1295257956.46, 1295258117.7,
  1295257956.46, 1295258117.7,
  1295258034.74, 1295258195.98,
  1295258034.74, 1295258195.98,
  1295258112.16, 1295258273.4,
  1295258112.16, 1295258273.4,
  1295258190.22, 1295258351.46,
  1295258190.22, 1295258351.46,
  1295258267.42, 1295258428.66,
  1295258267.42, 1295258428.66,
  1295258345.8, 1295258507.04,
  1295258345.8, 1295258507.04,
  1295258423.08, 1295258584.32,
  1295258423.08, 1295258584.32,
  1295258501.06, 1295258662.3,
  1295258501.06, 1295258662.3,
  1295258578.7, 1295258739.94,
  1295258578.7, 1295258739.94,
  1295258657.02, 1295258818.26,
  1295258657.02, 1295258818.26,
  1295258734.02, 1295258895.26,
  1295258734.02, 1295258895.26,
  1295258811.58, 1295258972.82,
  1295258811.58, 1295258972.82,
  1295258888.76, 1295259050,
  1295258888.76, 1295259050,
  1295258967.02, 1295259128.26,
  1295258967.02, 1295259128.26,
  1295259044.92, 1295259206.16,
  1295259044.92, 1295259206.16,
  1295259122.38, 1295259283.62,
  1295259122.38, 1295259283.62,
  1295259200.84, 1295259362.08,
  1295259200.84, 1295259362.08,
  1295259278.52, 1295259439.76,
  1295259278.52, 1295259439.76,
  1295259356.6, 1295259517.84,
  1295259356.6, 1295259517.84,
  1295259434.28, 1295259595.52,
  1295259434.28, 1295259595.52,
  1295259511.76, 1295259673,
  1295259511.76, 1295259673,
  1295259589.02, 1295259750.26,
  1295259589.02, 1295259750.26,
  1295259667.6, 1295259828.84,
  1295259667.6, 1295259828.84,
  1295259745.24, 1295259906.48,
  1295259745.24, 1295259906.48,
  1295259823.86, 1295259985.1,
  1295259823.86, 1295259985.1,
  1295259900.82, 1295260062.06,
  1295259900.82, 1295260062.06,
  1295259978.96, 1295260140.2,
  1295259978.96, 1295260140.2,
  1295260056.8, 1295260218.04,
  1295260056.8, 1295260218.04,
  1295260134.36, 1295260295.6,
  1295260134.36, 1295260295.6,
  1295260211.92, 1295260373.16,
  1295260211.92, 1295260373.16,
  1295260291.04, 1295260452.28,
  1295260291.04, 1295260452.28,
  1295260368, 1295260529.24,
  1295260368, 1295260529.24,
  1295260445.9, 1295260607.14,
  1295260445.9, 1295260607.14,
  1295260523.2, 1295260684.44,
  1295260523.2, 1295260684.44,
  1295260601.28, 1295260762.52,
  1295260601.28, 1295260762.52,
  1295260679.78, 1295260841.02,
  1295260679.78, 1295260841.02,
  1295260757.48, 1295260918.72,
  1295260757.48, 1295260918.72,
  1295260835.12, 1295260996.36,
  1295260835.12, 1295260996.36,
  1295260912.84, 1295261074.08,
  1295260912.84, 1295261074.08,
  1295260990.48, 1295261151.72,
  1295260990.48, 1295261151.72,
  1295261067.7, 1295261228.94,
  1295261067.7, 1295261228.94,
  1295261146.36, 1295261307.6,
  1295261146.36, 1295261307.6,
  1295261223.92, 1295261385.16,
  1295261223.92, 1295261385.16,
  1295261301.92, 1295261463.16,
  1295261301.92, 1295261463.16,
  1295261380.62, 1295261541.86,
  1295261380.62, 1295261541.86,
  1295261457.5, 1295261618.74,
  1295261457.5, 1295261618.74,
  1295261534.4, 1295261695.64,
  1295261534.4, 1295261695.64,
  1295261613.08, 1295261774.32,
  1295261613.08, 1295261774.32,
  1295261690.9, 1295261852.14,
  1295261690.9, 1295261852.14,
  1295261768.5, 1295261929.74,
  1295261768.5, 1295261929.74,
  1295261846.24, 1295262007.48,
  1295261846.24, 1295262007.48,
  1295261924.36, 1295262085.6,
  1295261924.36, 1295262085.6,
  1295262001.76, 1295262163,
  1295262001.76, 1295262163,
  1295262079.74, 1295262240.98,
  1295262079.74, 1295262240.98,
  1295262156.72, 1295262317.96,
  1295262156.72, 1295262317.96,
  1295262234.4, 1295262395.64,
  1295262234.4, 1295262395.64,
  1295262312.36, 1295262473.6,
  1295262312.36, 1295262473.6,
  1295262390.18, 1295262551.42,
  1295262390.18, 1295262551.42,
  1295262468.04, 1295262629.28,
  1295262468.04, 1295262629.28,
  1295262546.16, 1295262707.4,
  1295262546.16, 1295262707.4,
  1295262623.78, 1295262785.02,
  1295262623.78, 1295262785.02,
  1295262701.8, 1295262863.04,
  1295262701.8, 1295262863.04,
  1295262779.88, 1295262941.12,
  1295262779.88, 1295262941.12,
  1295262857.22, 1295263018.46,
  1295262857.22, 1295263018.46,
  1295262935.44, 1295263096.68,
  1295262935.44, 1295263096.68,
  1295263012.98, 1295263174.22,
  1295263012.98, 1295263174.22,
  1295263090.84, 1295263252.08,
  1295263090.84, 1295263252.08,
  1295263168.8, 1295263330.04,
  1295263168.8, 1295263330.04,
  1295263246.62, 1295263407.86,
  1295263246.62, 1295263407.86,
  1295263325.22, 1295263486.46,
  1295263325.22, 1295263486.46,
  1295263403.1, 1295263564.34,
  1295263403.1, 1295263564.34,
  1295263480.02, 1295263641.26,
  1295263480.02, 1295263641.26,
  1295263558.24, 1295263719.48,
  1295263558.24, 1295263719.48,
  1295263636.74, 1295263797.98,
  1295263636.74, 1295263797.98,
  1295263713.96, 1295263875.2,
  1295263713.96, 1295263875.2,
  1295263791.92, 1295263953.16,
  1295263791.92, 1295263953.16,
  1295263869, 1295264030.24,
  1295263869, 1295264030.24,
  1295263947.06, 1295264108.3,
  1295263947.06, 1295264108.3,
  1295264025.06, 1295264186.3,
  1295264025.06, 1295264186.3,
  1295264102.86, 1295264264.1,
  1295264102.86, 1295264264.1,
  1295264180.5, 1295264341.74,
  1295264180.5, 1295264341.74,
  1295264258.3, 1295264419.54,
  1295264258.3, 1295264419.54,
  1295264336.2, 1295264497.44,
  1295264336.2, 1295264497.44,
  1295264414.32, 1295264575.56,
  1295264414.32, 1295264575.56,
  1295264492.26, 1295264653.5,
  1295264492.26, 1295264653.5,
  1295264570.14, 1295264731.38,
  1295264570.14, 1295264731.38,
  1295264647.88, 1295264809.12,
  1295264647.88, 1295264809.12,
  1295264725.12, 1295264886.36,
  1295264725.12, 1295264886.36,
  1295264802.48, 1295264963.72,
  1295264802.48, 1295264963.72,
  1295264880.32, 1295265041.56,
  1295264880.32, 1295265041.56,
  1295264957.84, 1295265119.08,
  1295264957.84, 1295265119.08,
  1295265035.58, 1295265196.82,
  1295265035.58, 1295265196.82,
  1295265113.42, 1295265274.66,
  1295265113.42, 1295265274.66,
  1295265192.14, 1295265353.38,
  1295265192.14, 1295265353.38,
  1295265269.42, 1295265430.66,
  1295265269.42, 1295265430.66,
  1295265347.4, 1295265508.64,
  1295265347.4, 1295265508.64,
  1295265424.68, 1295265585.92,
  1295265424.68, 1295265585.92,
  1295265503.14, 1295265664.38,
  1295265503.14, 1295265664.38,
  1295265581.16, 1295265742.4,
  1295265581.16, 1295265742.4,
  1295265658.74, 1295265819.98,
  1295265658.74, 1295265819.98,
  1295265736.18, 1295265897.42,
  1295265736.18, 1295265897.42,
  1295265814.12, 1295265975.36,
  1295265814.12, 1295265975.36,
  1295265891.52, 1295266052.76,
  1295265891.52, 1295266052.76,
  1295265968.98, 1295266130.22,
  1295265968.98, 1295266130.22,
  1295266046.86, 1295266208.1,
  1295266046.86, 1295266208.1,
  1295266124.64, 1295266285.88,
  1295266124.64, 1295266285.88,
  1295266202.5, 1295266363.74,
  1295266202.5, 1295266363.74,
  1295266280.46, 1295266441.7,
  1295266280.46, 1295266441.7,
  1295266358.24, 1295266519.48,
  1295266358.24, 1295266519.48,
  1295266435.9, 1295266597.14,
  1295266435.9, 1295266597.14,
  1295266513.6, 1295266674.84,
  1295266513.6, 1295266674.84,
  1295266591.12, 1295266752.36,
  1295266591.12, 1295266752.36,
  1295266669.12, 1295266830.36,
  1295266669.12, 1295266830.36,
  1295266746.8, 1295266908.04,
  1295266746.8, 1295266908.04,
  1295266824.28, 1295266985.52,
  1295266824.28, 1295266985.52,
  1295266902.2, 1295267063.44,
  1295266902.2, 1295267063.44,
  1295266979.94, 1295267141.18,
  1295266979.94, 1295267141.18,
  1295267058.04, 1295267219.28,
  1295267058.04, 1295267219.28,
  1295267135.6, 1295267296.84,
  1295267135.6, 1295267296.84,
  1295267213.92, 1295267375.16,
  1295267213.92, 1295267375.16,
  1295267292.24, 1295267453.48,
  1295267292.24, 1295267453.48,
  1295267370.44, 1295267531.68,
  1295267370.44, 1295267531.68,
  1295267448.68, 1295267609.92,
  1295267448.68, 1295267609.92,
  1295267525.88, 1295267687.12,
  1295267525.88, 1295267687.12,
  1295267603.66, 1295267764.9,
  1295267603.66, 1295267764.9,
  1295267680.44, 1295267841.68,
  1295267680.44, 1295267841.68,
  1295267758, 1295267919.24,
  1295267758, 1295267919.24,
  1295267835.6, 1295267996.84,
  1295267835.6, 1295267996.84,
  1295267913.5, 1295268074.74,
  1295267913.5, 1295268074.74,
  1295267991.06, 1295268152.3,
  1295267991.06, 1295268152.3,
  1295268068.32, 1295268229.56,
  1295268068.32, 1295268229.56,
  1295268145.9, 1295268307.14,
  1295268145.9, 1295268307.14,
  1295268227.5, 1295268388.74,
  1295268227.5, 1295268388.74,
  1295268303.62, 1295268464.86,
  1295268303.62, 1295268464.86,
  1295268381.4, 1295268542.64,
  1295268381.4, 1295268542.64,
  1295268458.88, 1295268620.12,
  1295268458.88, 1295268620.12,
  1295268537.6, 1295268698.84,
  1295268537.6, 1295268698.84,
  1295268615.46, 1295268776.7,
  1295268615.46, 1295268776.7,
  1295268693.94, 1295268855.18,
  1295268693.94, 1295268855.18,
  1295268770.9, 1295268932.14,
  1295268770.9, 1295268932.14,
  1295268849.26, 1295269010.5,
  1295268849.26, 1295269010.5,
  1295268927.26, 1295269088.5,
  1295268927.26, 1295269088.5,
  1295269005.34, 1295269166.58,
  1295269005.34, 1295269166.58,
  1295269082.84, 1295269244.08,
  1295269082.84, 1295269244.08,
  1295269162.26, 1295269323.5,
  1295269162.26, 1295269323.5,
  1295269239.44, 1295269400.68,
  1295269239.44, 1295269400.68,
  1295269317.66, 1295269478.9,
  1295269317.66, 1295269478.9,
  1295269394.9, 1295269556.14,
  1295269394.9, 1295269556.14,
  1295269473.16, 1295269634.4,
  1295269473.16, 1295269634.4,
  1295269551.14, 1295269712.38,
  1295269551.14, 1295269712.38,
  1295269628.06, 1295269789.3,
  1295269628.06, 1295269789.3,
  1295269705.52, 1295269866.76,
  1295269705.52, 1295269866.76,
  1295269782.98, 1295269944.22,
  1295269782.98, 1295269944.22,
  1295269859.2, 1295270020.44,
  1295269859.2, 1295270020.44,
  1295269936.62, 1295270097.86,
  1295269936.62, 1295270097.86,
  1295270013.82, 1295270175.06,
  1295270013.82, 1295270175.06,
  1295270091.68, 1295270252.92,
  1295270091.68, 1295270252.92,
  1295270170.4, 1295270331.64,
  1295270170.4, 1295270331.64,
  1295270249, 1295270410.24,
  1295270249, 1295270410.24,
  1295270326.88, 1295270488.12,
  1295270326.88, 1295270488.12,
  1295270407.82, 1295270569.06,
  1295270407.82, 1295270569.06,
  1295270483.64, 1295270644.88,
  1295270483.64, 1295270644.88,
  1295270561.08, 1295270722.32,
  1295270561.08, 1295270722.32,
  1295270640.52, 1295270801.76,
  1295270640.52, 1295270801.76,
  1295270717.86, 1295270879.1,
  1295270717.86, 1295270879.1,
  1295270794.58, 1295270955.82,
  1295270794.58, 1295270955.82,
  1295270872.2, 1295271033.44,
  1295270872.2, 1295271033.44,
  1295270949.68, 1295271110.92,
  1295270949.68, 1295271110.92,
  1295271028.02, 1295271189.26,
  1295271028.02, 1295271189.26,
  1295271105.4, 1295271266.64,
  1295271105.4, 1295271266.64,
  1295271182.16, 1295271343.4,
  1295271182.16, 1295271343.4,
  1295271259.22, 1295271420.46,
  1295271259.22, 1295271420.46,
  1295271336.06, 1295271497.3,
  1295271336.06, 1295271497.3,
  1295271413.72, 1295271574.96,
  1295271413.72, 1295271574.96,
  1295271492.34, 1295271653.58,
  1295271492.34, 1295271653.58,
  1295271570.1, 1295271731.34,
  1295271570.1, 1295271731.34,
  1295271645.98, 1295271807.22,
  1295271645.98, 1295271807.22,
  1295271723.22, 1295271884.46,
  1295271723.22, 1295271884.46,
  1295271801.3, 1295271962.54,
  1295271801.3, 1295271962.54,
  1295271878.84, 1295272040.08,
  1295271878.84, 1295272040.08,
  1295271956.32, 1295272117.56,
  1295271956.32, 1295272117.56,
  1295272034.28, 1295272195.52,
  1295272034.28, 1295272195.52,
  1295272113.14, 1295272274.38,
  1295272113.14, 1295272274.38,
  1295272192.04, 1295272353.28,
  1295272192.04, 1295272353.28,
  1295272270.38, 1295272431.62,
  1295272270.38, 1295272431.62,
  1295272348.72, 1295272509.96,
  1295272348.72, 1295272509.96,
  1295272427.14, 1295272588.38,
  1295272427.14, 1295272588.38,
  1295272504.68, 1295272665.92,
  1295272504.68, 1295272665.92,
  1295272582.12, 1295272743.36,
  1295272582.12, 1295272743.36,
  1295272658.58, 1295272819.82,
  1295272658.58, 1295272819.82,
  1295272735.68, 1295272896.92,
  1295272735.68, 1295272896.92,
  1295272811.78, 1295272973.02,
  1295272811.78, 1295272973.02,
  1295272889.2, 1295273050.44,
  1295272889.2, 1295273050.44,
  1295272966.98, 1295273128.22,
  1295272966.98, 1295273128.22,
  1295273045.32, 1295273206.56,
  1295273045.32, 1295273206.56,
  1295273125.26, 1295273286.5,
  1295273125.26, 1295273286.5,
  1295273203.52, 1295273364.76,
  1295273203.52, 1295273364.76,
  1295273281.22, 1295273442.46,
  1295273281.22, 1295273442.46,
  1295273357.82, 1295273519.06,
  1295273357.82, 1295273519.06,
  1295273433.76, 1295273595,
  1295273433.76, 1295273595,
  1295273509.26, 1295273670.5,
  1295273509.26, 1295273670.5,
  1295273585.88, 1295273747.12,
  1295273585.88, 1295273747.12,
  1295273662.04, 1295273823.28,
  1295273662.04, 1295273823.28,
  1295273740.24, 1295273901.48,
  1295273740.24, 1295273901.48,
  1295273818.64, 1295273979.88,
  1295273818.64, 1295273979.88,
  1295273897.84, 1295274059.08,
  1295273897.84, 1295274059.08,
  1295273976, 1295274137.24,
  1295273976, 1295274137.24,
  1295274052.64, 1295274213.88,
  1295274052.64, 1295274213.88,
  1295274130.46, 1295274291.7,
  1295274130.46, 1295274291.7,
  1295274208.16, 1295274369.4,
  1295274208.16, 1295274369.4,
  1295274287.84, 1295274449.08,
  1295274287.84, 1295274449.08,
  1295274366.88, 1295274528.12,
  1295274366.88, 1295274528.12,
  1295274445.98, 1295274607.22,
  1295274445.98, 1295274607.22,
  1295274522.8, 1295274684.04,
  1295274522.8, 1295274684.04,
  1295274598.86, 1295274760.1,
  1295274598.86, 1295274760.1,
  1295274675.76, 1295274837,
  1295274675.76, 1295274837,
  1295274754.62, 1295274915.86,
  1295274754.62, 1295274915.86,
  1295274832.12, 1295274993.36,
  1295274832.12, 1295274993.36,
  1295274909.32, 1295275070.56,
  1295274909.32, 1295275070.56,
  1295274988.4, 1295275149.64,
  1295274988.4, 1295275149.64,
  1295275066.28, 1295275227.52,
  1295275066.28, 1295275227.52,
  1295275142.64, 1295275303.88,
  1295275142.64, 1295275303.88,
  1295275220.48, 1295275381.72,
  1295275220.48, 1295275381.72,
  1295275298.4, 1295275459.64,
  1295275298.4, 1295275459.64,
  1295275376.48, 1295275537.72,
  1295275376.48, 1295275537.72,
  1295275455.38, 1295275616.62,
  1295275455.38, 1295275616.62,
  1295275534.7, 1295275695.94,
  1295275534.7, 1295275695.94,
  1295275613.3, 1295275774.54,
  1295275613.3, 1295275774.54,
  1295275690.46, 1295275851.7,
  1295275690.46, 1295275851.7,
  1295275768.6, 1295275929.84,
  1295275768.6, 1295275929.84,
  1295275846.2, 1295276007.44,
  1295275846.2, 1295276007.44,
  1295275921.96, 1295276083.2,
  1295275921.96, 1295276083.2,
  1295276000, 1295276161.24,
  1295276000, 1295276161.24,
  1295276076.9, 1295276238.14,
  1295276076.9, 1295276238.14,
  1295276154.22, 1295276315.46,
  1295276154.22, 1295276315.46,
  1295276232.36, 1295276393.6,
  1295276232.36, 1295276393.6,
  1295276309.94, 1295276471.18,
  1295276309.94, 1295276471.18,
  1295276386.98, 1295276548.22,
  1295276386.98, 1295276548.22,
  1295276464.44, 1295276625.68,
  1295276464.44, 1295276625.68,
  1295276542.24, 1295276703.48,
  1295276542.24, 1295276703.48,
  1295276620, 1295276781.24,
  1295276620, 1295276781.24,
  1295276697.98, 1295276859.22,
  1295276697.98, 1295276859.22,
  1295276774.92, 1295276936.16,
  1295276774.92, 1295276936.16,
  1295276853.78, 1295277015.02,
  1295276853.78, 1295277015.02,
  1295276931.54, 1295277092.78,
  1295276931.54, 1295277092.78,
  1295277009.98, 1295277171.22,
  1295277009.98, 1295277171.22,
  1295277087.32, 1295277248.56,
  1295277087.32, 1295277248.56,
  1295277166.1, 1295277327.34,
  1295277166.1, 1295277327.34,
  1295277243.38, 1295277404.62,
  1295277243.38, 1295277404.62,
  1295277321.7, 1295277482.94,
  1295277321.7, 1295277482.94,
  1295277399.58, 1295277560.82,
  1295277399.58, 1295277560.82,
  1295277477.02, 1295277638.26,
  1295277477.02, 1295277638.26,
  1295277555.9, 1295277717.14,
  1295277555.9, 1295277717.14,
  1295277634.92, 1295277796.16,
  1295277634.92, 1295277796.16,
  1295277712.96, 1295277874.2,
  1295277712.96, 1295277874.2,
  1295277791.18, 1295277952.42,
  1295277791.18, 1295277952.42,
  1295277868.98, 1295278030.22,
  1295277868.98, 1295278030.22,
  1295277946.72, 1295278107.96,
  1295277946.72, 1295278107.96,
  1295278024.02, 1295278185.26,
  1295278024.02, 1295278185.26 ;

 emf =
  3.998894e-014, 3.666264e-015, -3.832919e-011, 5.610733e-012,
  3.195066e-014, 4.172533e-015, -6.178277e-011, 6.316628e-011,
  3.569003e-014, 4.605785e-015, 5.446329e-011, 6.15795e-011,
  2.818398e-014, 2.086935e-015, 3.866479e-011, 1.431981e-010,
  1.056961e-013, -7.815512e-015, 1.222013e-012, 1.027887e-011,
  1.488394e-014, 3.87379e-015, -1.482599e-011, 7.083661e-011,
  1.384893e-013, -1.296095e-014, 6.092587e-011, 8.197641e-011,
  9.5958e-014, -4.702634e-015, -5.183726e-011, 5.312005e-011,
  4.924692e-014, 2.658534e-015, 6.063121e-011, 9.78786e-011,
  3.931066e-014, 2.25092e-015, -9.702908e-012, 8.48524e-011,
  3.534706e-014, 4.197324e-015, -2.391802e-011, 7.155844e-012,
  3.411273e-014, 3.812066e-015, 2.167501e-011, 1.02676e-010,
  -2.260401e-014, 1.386701e-014, -9.781797e-011, -2.127638e-011,
  -3.477418e-015, 1.090597e-014, -2.183201e-011, 4.882823e-011,
  3.803661e-014, 6.481471e-015, -1.619536e-011, 5.280348e-011,
  3.935748e-014, 6.639484e-015, -5.491792e-011, 5.865584e-011,
  4.272083e-014, 5.562069e-015, -9.96796e-011, -2.115693e-012,
  3.267036e-014, 7.655299e-015, 5.73925e-012, 1.022014e-010,
  4.027253e-014, 2.360733e-014, -1.440128e-011, 2.476691e-011,
  2.061508e-015, -8.779018e-015, -2.287384e-011, 7.137393e-011,
  2.014655e-014, 1.124736e-014, 4.473687e-011, 8.46681e-011,
  -2.721147e-014, 1.771517e-014, 3.480146e-011, 1.540384e-010,
  3.850938e-014, 9.009075e-015, 8.429269e-012, 6.508991e-011,
  3.363913e-014, 9.284664e-015, 7.316522e-012, 8.748498e-011,
  5.493917e-014, 6.552838e-015, -1.055587e-011, 6.286593e-011,
  1.745732e-013, -1.113551e-014, 5.10395e-012, 1.113264e-010,
  4.343299e-014, 7.540757e-015, 9.042301e-012, 6.662872e-011,
  7.030977e-014, 4.979648e-015, -3.440625e-011, 1.001467e-010,
  4.075285e-014, 8.474814e-015, 2.658599e-011, 1.092462e-010,
  5.603652e-014, 7.96622e-015, -1.174512e-011, 1.387049e-010,
  3.794294e-014, 8.360366e-015, 6.926681e-013, 5.304464e-011,
  5.312591e-014, 1.113044e-014, -5.000839e-011, 1.334687e-010,
  1.78385e-014, 1.236325e-014, 5.911281e-011, 9.069788e-011,
  4.507131e-014, 1.069153e-014, 4.405889e-011, 2.038982e-010,
  4.796382e-014, 8.569562e-015, 5.189565e-012, 5.701981e-011,
  6.284049e-014, 7.546644e-015, -1.313614e-010, 5.415331e-011,
  4.181539e-014, 7.380873e-015, -8.856516e-012, 5.495776e-011,
  4.963581e-014, 1.116246e-014, -1.313864e-011, 7.319939e-011,
  4.148092e-014, 7.755222e-015, 8.821689e-012, 9.066085e-011,
  5.843766e-014, 8.519025e-015, -6.505431e-011, 7.720252e-011,
  4.144276e-014, 7.372985e-015, 4.347827e-011, 7.915844e-011,
  6.328001e-014, 8.805387e-015, -2.701375e-011, 1.185186e-010,
  4.314192e-014, 7.714663e-015, 5.186618e-011, 9.2276e-011,
  6.18024e-014, 7.423457e-015, 4.227023e-011, 1.327712e-010,
  4.852459e-014, 5.70255e-015, -2.734317e-011, 4.884639e-011,
  6.832952e-014, 4.939e-015, -3.221265e-013, 1.247416e-010,
  6.371955e-014, 2.598917e-015, 6.333014e-012, 1.071079e-010,
  6.257715e-014, 2.70354e-015, -4.599341e-011, 7.971319e-011,
  6.376755e-014, 8.840389e-015, -2.206689e-011, 1.173039e-010,
  7.91057e-014, 2.319111e-015, -2.600844e-011, 1.434725e-010,
  5.968542e-014, 5.759884e-015, -1.334477e-011, 8.661893e-011,
  1.027859e-013, -7.757355e-016, -1.060898e-010, 8.729117e-011,
  5.484701e-014, 2.17714e-015, -6.068606e-011, 4.805886e-011,
  8.978426e-014, 1.606699e-015, -4.467667e-011, 1.421618e-010,
  1.085269e-013, -5.948546e-015, 1.847706e-011, 8.845871e-011,
  1.144045e-013, -4.626515e-015, 7.489987e-012, 1.411885e-010,
  3.525782e-014, 4.898896e-015, 2.794739e-011, 7.315485e-011,
  9.459969e-014, -2.838907e-015, -1.986164e-011, 1.471536e-010,
  2.086549e-014, 5.798452e-015, 9.813881e-011, 1.019704e-010,
  8.915991e-014, -2.468415e-015, 4.38378e-011, 2.236594e-010,
  4.462136e-014, 3.126387e-015, 9.264657e-011, 1.325966e-010,
  1.080646e-013, -4.994983e-015, -2.995057e-011, 1.12086e-010,
  5.469643e-014, 3.317888e-015, 5.357495e-011, 2.141805e-010,
  1.149698e-013, -4.627193e-015, 1.205796e-011, 1.443483e-010,
  4.903993e-014, 4.860363e-015, 2.511567e-011, 1.249269e-010,
  1.212784e-013, -3.172012e-015, 6.477968e-011, 2.218069e-010,
  6.015636e-014, 4.517225e-015, -5.657443e-011, 5.113867e-011,
  1.178877e-013, -9.65987e-017, 1.088832e-010, 2.58331e-010,
  5.695418e-014, 4.072198e-015, -1.038947e-010, 1.067605e-011,
  1.367265e-013, -2.338925e-015, -3.757552e-011, 1.492152e-010,
  2.975386e-014, 1.023849e-014, -1.371879e-011, 1.002743e-010,
  1.202196e-013, -6.711158e-016, 1.165224e-010, 2.635378e-010,
  5.002293e-014, 5.410701e-015, -4.153384e-011, 1.071428e-010,
  1.474862e-013, -6.858214e-015, 4.91177e-011, 2.315601e-010,
  4.48294e-014, 5.587306e-015, 7.902304e-011, 1.293871e-010,
  1.664295e-013, -8.062159e-015, 3.045051e-011, 2.299912e-010,
  6.88182e-014, 6.041396e-015, -7.379244e-011, 8.25841e-011,
  1.621371e-013, 9.058419e-017, 5.69475e-011, 2.066156e-010,
  5.97966e-014, 1.072393e-014, -1.969745e-011, 1.105246e-010,
  1.566767e-013, 1.11951e-014, -3.864993e-011, 1.950409e-010,
  5.306596e-014, 1.741614e-014, 4.663269e-011, 1.919123e-010,
  1.264587e-013, 2.223411e-014, -1.397551e-011, 2.531471e-010,
  6.396499e-014, 1.743255e-014, 1.611939e-011, 1.358629e-010,
  1.876453e-013, 1.668778e-014, 4.930548e-011, 2.732108e-010,
  6.524929e-014, 1.842837e-014, -1.903972e-011, 1.361813e-010,
  2.061349e-013, 2.031054e-014, 5.494784e-011, 2.694387e-010,
  6.760045e-014, 2.178348e-014, -8.434566e-011, 9.738089e-011,
  2.210743e-013, 2.325281e-014, -9.39556e-011, 1.948941e-010,
  1.143572e-013, 1.663853e-014, -4.006395e-011, 1.196714e-010,
  1.694375e-013, 3.579745e-014, 5.671724e-013, 2.341277e-010,
  7.332416e-014, 2.860226e-014, -8.671303e-011, 9.792366e-011,
  2.439992e-013, 3.397798e-014, 2.755103e-012, 2.490151e-010,
  7.099309e-014, 3.254774e-014, -2.519199e-011, 1.614339e-010,
  2.631288e-013, 3.97723e-014, -8.82932e-011, 2.007867e-010,
  6.616012e-014, 4.012651e-014, 7.661193e-011, 2.399545e-010,
  2.734946e-013, 5.269076e-014, -7.661444e-011, 2.253304e-010,
  8.107043e-014, 3.491714e-014, 3.672378e-012, 2.519519e-010,
  2.952432e-013, 6.353797e-014, -6.154947e-011, 3.082731e-010,
  9.077164e-014, 5.292472e-014, -3.701624e-011, 2.063894e-010,
  3.071577e-013, 7.288143e-014, -7.157414e-011, 2.717141e-010,
  9.919731e-014, 5.442466e-014, -9.775269e-011, 1.964197e-010,
  3.39414e-013, 7.180376e-014, -1.075051e-010, 2.625774e-010,
  1.143586e-013, 5.090538e-014, -1.363466e-010, 1.576385e-010,
  3.449598e-013, 6.589836e-014, -7.1315e-012, 2.961011e-010,
  1.644774e-013, 4.128277e-014, -9.143942e-011, 2.06694e-010,
  3.697594e-013, 6.003961e-014, -4.199951e-011, 3.204172e-010,
  1.42713e-013, 4.572251e-014, 1.844291e-011, 3.233772e-010,
  4.021254e-013, 5.407877e-014, -1.340349e-010, 2.838464e-010,
  1.133023e-013, 4.933059e-014, -3.881917e-011, 2.028962e-010,
  4.242901e-013, 5.018703e-014, -5.053915e-011, 3.277335e-010,
  1.335351e-013, 4.213637e-014, -3.910536e-011, 2.508626e-010,
  4.702773e-013, 3.650286e-014, -1.093602e-010, 2.807767e-010,
  1.474325e-013, 3.914802e-014, 3.755071e-011, 2.860241e-010,
  4.968828e-013, 2.970184e-014, -1.409247e-011, 3.450666e-010,
  1.958192e-013, 3.184401e-014, -6.383041e-011, 2.311244e-010,
  5.561586e-013, 2.005566e-014, -7.173694e-011, 2.958996e-010,
  1.620591e-013, 3.398552e-014, 5.548414e-011, 3.432014e-010,
  5.615999e-013, 1.565429e-014, 4.264351e-013, 3.510968e-010,
  1.780035e-013, 2.858219e-014, -2.269253e-011, 2.971354e-010,
  5.907461e-013, 7.213048e-015, -5.099323e-011, 3.661389e-010,
  1.86808e-013, 2.095194e-014, 7.411818e-011, 3.433629e-010,
  6.296349e-013, -6.812715e-015, -4.826817e-011, 3.607389e-010,
  2.174462e-013, 1.496837e-014, -4.797008e-011, 3.01685e-010,
  6.579571e-013, -1.311723e-014, 1.171284e-010, 4.475874e-010,
  2.385979e-013, 1.521519e-014, -6.332258e-011, 3.125792e-010,
  7.172638e-013, -1.506445e-014, -4.073127e-012, 3.855282e-010,
  2.444625e-013, 1.821154e-014, 6.439671e-011, 4.257126e-010,
  7.654672e-013, -1.598573e-014, 8.899459e-012, 4.159478e-010,
  2.798993e-013, 1.490814e-014, -1.970427e-011, 3.987616e-010,
  8.231576e-013, -1.970126e-014, -1.650517e-011, 4.147532e-010,
  3.009943e-013, 1.42901e-014, 1.192794e-011, 4.14879e-010,
  8.726734e-013, -2.259292e-014, -8.287046e-011, 4.114601e-010,
  3.255811e-013, 1.382673e-014, 3.859903e-011, 4.190568e-010,
  9.298197e-013, -2.512693e-014, -1.068259e-011, 4.232038e-010,
  3.605045e-013, 1.500846e-014, 3.197557e-011, 4.631037e-010,
  1.001449e-012, -2.436326e-014, 6.939014e-011, 5.286195e-010,
  4.046795e-013, 1.764347e-014, -4.304542e-011, 4.417055e-010,
  1.077086e-012, -2.263496e-014, 4.229506e-011, 4.868854e-010,
  4.073938e-013, 2.701859e-014, 6.298903e-012, 5.044485e-010,
  1.195468e-012, -2.438872e-014, -2.994476e-011, 4.717861e-010,
  4.731344e-013, 2.904631e-014, 8.540385e-011, 5.931697e-010,
  1.235133e-012, -2.030706e-014, 5.982202e-011, 5.235044e-010,
  5.283818e-013, 2.974642e-014, -8.052647e-011, 5.17308e-010,
  1.305429e-012, -1.662269e-014, 9.37426e-011, 5.618266e-010,
  5.923931e-013, 2.085115e-014, -5.496701e-011, 5.475784e-010,
  1.397496e-012, -2.458334e-014, 4.379738e-011, 5.890524e-010,
  6.713913e-013, 1.096679e-014, -6.405688e-011, 5.632768e-010,
  1.46831e-012, -2.879914e-014, 2.981125e-011, 6.000191e-010,
  7.492145e-013, 1.979216e-014, -2.807932e-011, 6.134624e-010,
  1.559645e-012, -2.138411e-014, 5.96244e-011, 6.305561e-010,
  7.997985e-013, 4.885631e-014, -1.061028e-010, 6.335193e-010,
  1.704624e-012, -8.745427e-015, 3.401893e-011, 6.400375e-010,
  8.761719e-013, 6.721099e-014, -2.680588e-011, 7.004021e-010,
  1.829774e-012, 2.813869e-015, 1.218789e-011, 6.577775e-010,
  9.746342e-013, 5.551432e-014, -1.206983e-010, 6.436963e-010,
  1.955457e-012, -8.662245e-015, 4.304677e-011, 6.64883e-010,
  1.086237e-012, 1.852508e-014, -4.990382e-013, 8.351515e-010,
  2.083978e-012, -3.957719e-014, 5.409697e-011, 6.595594e-010,
  1.200913e-012, -6.791743e-015, 6.768364e-011, 8.666731e-010,
  2.230128e-012, -6.238905e-014, -2.120504e-011, 6.757664e-010,
  1.331102e-012, 5.955789e-016, -3.40275e-011, 8.242501e-010,
  2.392333e-012, -6.112392e-014, 9.858389e-012, 6.403237e-010,
  1.484055e-012, 3.232004e-014, 6.728177e-012, 9.003278e-010,
  2.573251e-012, -4.214155e-014, 4.298101e-011, 7.12934e-010,
  1.654243e-012, 6.017798e-014, -1.410028e-010, 8.525954e-010,
  2.745747e-012, -2.420716e-014, 2.33205e-011, 7.426087e-010,
  1.834342e-012, 4.071244e-014, 4.606196e-011, 1.051232e-009,
  2.965436e-012, -4.610637e-014, 5.250218e-013, 7.189336e-010,
  2.039781e-012, 4.116703e-015, 4.078265e-011, 1.10452e-009,
  3.181324e-012, -7.223659e-014, 2.600143e-011, 7.552728e-010,
  2.287648e-012, -1.492986e-014, 5.883907e-011, 1.150475e-009,
  3.417506e-012, -8.893427e-014, -1.945529e-011, 7.648376e-010,
  2.600107e-012, -4.064098e-014, 2.823062e-011, 1.167034e-009,
  3.733496e-012, -1.112152e-013, 3.263858e-011, 7.394961e-010,
  2.867556e-012, -4.385139e-014, 1.485107e-010, 1.316736e-009,
  3.965475e-012, -1.097186e-013, 5.356291e-012, 8.149033e-010,
  3.193236e-012, -7.840477e-014, 4.084754e-011, 1.266686e-009,
  4.267701e-012, -1.293348e-013, 5.852911e-011, 8.164102e-010,
  3.57833e-012, -1.3071e-013, 6.609807e-011, 1.339835e-009,
  4.587579e-012, -1.544059e-013, 4.254471e-011, 8.121921e-010,
  4.015796e-012, -1.84732e-013, 2.193873e-010, 1.479376e-009,
  4.997843e-012, -1.913559e-013, 6.664739e-011, 8.580219e-010,
  4.49345e-012, -1.524721e-013, 6.003217e-011, 1.478682e-009,
  5.349567e-012, -1.757074e-013, 1.43097e-010, 8.920651e-010,
  5.034689e-012, -9.583424e-014, 1.341529e-010, 1.599952e-009,
  5.718433e-012, -1.500075e-013, 1.000245e-010, 8.866137e-010,
  5.670228e-012, -7.210016e-014, 4.319868e-011, 1.607671e-009,
  6.165235e-012, -1.445528e-013, 7.591577e-011, 8.756919e-010,
  6.373431e-012, -1.146899e-013, -5.818797e-011, 1.598267e-009,
  6.656576e-012, -1.63808e-013, 7.208546e-011, 8.343426e-010,
  7.166487e-012, -1.805377e-013, 4.109178e-011, 1.692094e-009,
  7.178424e-012, -1.952623e-013, 3.515818e-011, 7.526631e-010,
  8.056735e-012, -1.932671e-013, 5.711214e-011, 1.781308e-009,
  7.736258e-012, -2.057282e-013, 9.313805e-011, 7.860407e-010,
  9.087873e-012, -1.495265e-013, -4.836106e-011, 1.80096e-009,
  8.341664e-012, -1.987784e-013, 3.520655e-011, 7.470655e-010,
  1.02586e-011, -1.245299e-013, -7.914259e-011, 1.817946e-009,
  9.008456e-012, -2.002523e-013, 5.966782e-012, 6.983574e-010,
  1.158896e-011, -1.482758e-013, -9.903994e-012, 1.867336e-009,
  9.725562e-012, -2.139219e-013, 1.079799e-010, 7.352541e-010,
  1.314197e-011, -5.104395e-014, 1.44859e-011, 1.973878e-009,
  1.051998e-011, -1.965649e-013, 4.876561e-011, 6.454033e-010,
  1.490275e-011, 5.926543e-014, 8.070535e-012, 1.994604e-009,
  1.138204e-011, -1.785233e-013, 2.904415e-011, 6.014046e-010,
  1.693885e-011, 6.253588e-014, -4.410578e-011, 1.936161e-009,
  1.231474e-011, -1.819795e-013, 3.813936e-011, 5.070435e-010,
  1.933417e-011, -1.504601e-014, -9.228766e-011, 1.8278e-009,
  1.336939e-011, -1.96587e-013, 2.914947e-011, 4.139067e-010,
  2.209433e-011, -4.898897e-014, -5.497278e-011, 1.759878e-009,
  1.452877e-011, -2.002088e-013, 4.028967e-011, 3.094304e-010,
  2.529914e-011, -6.086172e-014, -4.40826e-011, 1.664332e-009,
  1.581107e-011, -1.955021e-013, 4.397907e-011, 2.410104e-010,
  2.917679e-011, -8.815259e-014, -3.494891e-011, 1.451229e-009,
  1.72326e-011, -1.887734e-013, 8.066374e-012, 4.374201e-011,
  3.367526e-011, -2.890879e-013, 9.089847e-011, 1.245135e-009,
  1.881194e-011, -1.987836e-013, -5.683969e-011, -1.396621e-010,
  3.901361e-011, -6.099126e-013, 2.279746e-010, 9.518826e-010,
  2.05815e-011, -2.211264e-013, 4.999552e-011, -3.459286e-010,
  4.529358e-011, -6.383197e-013, 6.445611e-011, 3.621111e-010,
  2.252297e-011, -2.111627e-013, -2.802781e-011, -5.959634e-010,
  5.287569e-011, -6.602245e-013, 1.06814e-010, -2.827731e-010,
  2.470666e-011, -2.026155e-013, 1.196838e-010, -7.548492e-010,
  6.194947e-011, -9.167368e-013, 1.304129e-010, -1.144347e-009,
  2.712639e-011, -2.006515e-013, -1.69012e-012, -1.199088e-009,
  7.302991e-011, -1.440688e-012, 3.000325e-010, -2.24705e-009,
  2.98739e-011, -2.059548e-013, 4.82961e-011, -1.597324e-009,
  8.648093e-011, -1.99609e-012, 3.972054e-010, -3.713911e-009,
  3.293388e-011, -2.070618e-013, 4.013044e-011, -2.035571e-009,
  1.03235e-010, -2.664226e-012, 5.73978e-010, -5.660509e-009,
  3.645404e-011, -1.837815e-013, 1.374675e-010, -2.523257e-009,
  1.241765e-010, -3.209897e-012, 5.333051e-010, -8.395246e-009,
  4.048463e-011, -1.289702e-013, 1.525999e-010, -3.174084e-009,
  1.505845e-010, -4.661834e-012, 6.954676e-010, -1.191556e-008,
  4.515475e-011, -8.326866e-014, 2.17597e-010, -3.899831e-009,
  1.841216e-010, -6.569829e-012, 1.026981e-009, -1.647447e-008,
  5.045509e-011, -1.58513e-014, 1.763677e-010, -4.843327e-009,
  2.255332e-010, -8.075629e-012, 9.132479e-010, -2.277956e-008,
  5.52679e-011, -1.320341e-013, 1.461155e-010, -5.9469e-009,
  2.853667e-010, -9.644732e-012, 1.029214e-009, -3.130735e-008,
  6.411138e-011, -1.819305e-013, 1.713031e-010, -7.238437e-009,
  3.651645e-010, -1.349119e-011, 1.334645e-009, -4.338053e-008,
  7.132747e-011, 3.17681e-013, 1.705177e-010, -8.932171e-009,
  4.778863e-010, -1.710361e-011, 1.584072e-009, -6.06399e-008,
  8.219395e-011, 4.849168e-013, 1.770224e-010, -1.097269e-008,
  6.40912e-010, -2.12603e-011, 1.682825e-009, -8.574164e-008,
  9.547965e-011, 6.170523e-013, 2.692879e-010, -1.346629e-008,
  8.934399e-010, -2.615608e-011, 2.096961e-009, -1.245796e-007,
  1.130124e-010, 8.792986e-013, 2.496057e-010, -1.679346e-008,
  1.304934e-009, -3.132112e-011, 2.830963e-009, -1.874587e-007,
  1.368648e-010, 1.478101e-012, 3.611617e-010, -2.151225e-008,
  2.021807e-009, -5.014502e-011, 6.442305e-009, -2.983307e-007,
  1.705122e-010, 2.012604e-012, 7.141501e-010, -2.820556e-008,
  3.280424e-009, -1.002881e-010, 1.631354e-008, -5.180945e-007,
  2.181562e-010, 2.909812e-012, 9.928643e-010, -3.838984e-008,
  4.48078e-009, -2.51218e-010, 4.129815e-008, -1.028792e-006,
  2.26285e-010, 2.69088e-012, 3.099903e-009, -5.782065e-008,
  -6.253438e-010, -5.492963e-010, 1.109757e-007, -2.210836e-006,
  3.203684e-011, 3.914748e-012, 5.398007e-009, -8.797555e-008,
  -1.036915e-008, -5.784933e-010, 1.718782e-007, -3.604822e-006,
  1.197321e-010, 1.191918e-011, 5.201999e-009, -9.132734e-008,
  -1.236542e-008, -5.802294e-010, 1.698424e-007, -4.019754e-006,
  2.378864e-010, 3.788699e-012, 2.965555e-009, -7.444786e-008,
  -9.379898e-009, -1.002209e-009, 1.155536e-007, -3.394451e-006,
  3.811397e-010, -9.481485e-012, 1.173156e-009, -4.698989e-008,
  7.972753e-010, -1.081183e-009, 5.009056e-008, -1.967655e-006,
  4.251949e-010, 9.451875e-012, 7.107883e-010, -2.563749e-008,
  4.526288e-009, -4.300678e-010, 1.927581e-008, -9.146281e-007,
  2.10339e-010, 1.195784e-011, 8.216279e-010, -2.651936e-008,
  3.122668e-009, -8.718772e-011, 6.941836e-009, -4.7291e-007,
  1.519584e-010, 5.087983e-012, 4.215275e-010, -2.506691e-008,
  1.92335e-009, -1.446545e-011, 2.057822e-009, -2.789425e-007,
  1.312039e-010, 8.208693e-013, 1.463572e-010, -2.113792e-008,
  1.248086e-009, -1.947063e-011, 1.123394e-009, -1.781409e-007,
  1.140032e-010, -6.458517e-014, 1.011189e-010, -1.753064e-008,
  8.632313e-010, -2.59342e-011, 1.316849e-009, -1.204366e-007,
  9.897056e-011, -2.88605e-013, 1.455723e-010, -1.455245e-008,
  6.262186e-010, -2.933393e-011, 2.140836e-009, -8.452137e-008,
  8.657906e-011, -8.449877e-014, 2.980173e-010, -1.207951e-008,
  4.698216e-010, -2.360977e-011, 2.239364e-009, -6.072047e-008,
  7.616877e-011, 1.200908e-013, 4.448561e-010, -9.901052e-009,
  3.628603e-010, -1.506136e-011, 1.809426e-009, -4.452356e-008,
  6.742185e-011, 1.584247e-013, 2.186201e-010, -8.356928e-009,
  2.861511e-010, -8.369138e-012, 1.451101e-009, -3.292104e-008,
  6.004258e-011, 1.509428e-013, 3.644424e-010, -6.899415e-009,
  2.291601e-010, -7.261709e-012, 1.300794e-009, -2.452768e-008,
  5.375448e-011, 8.555213e-014, 2.293877e-010, -5.860226e-009,
  1.87428e-010, -5.513195e-012, 1.381127e-009, -1.828411e-008,
  4.939955e-011, 1.780041e-013, 1.442511e-010, -4.846611e-009,
  1.540981e-010, -4.937007e-012, 1.327598e-009, -1.368425e-008,
  4.447637e-011, 1.999194e-013, 2.757216e-010, -3.972584e-009,
  1.278629e-010, -3.532617e-012, 1.126683e-009, -1.00613e-008,
  4.015249e-011, 2.554925e-013, 2.126529e-010, -3.330731e-009,
  1.068099e-010, -1.535682e-012, 8.049805e-010, -7.308379e-009,
  3.631209e-011, 3.251909e-013, 1.677839e-010, -2.656903e-009,
  8.981965e-011, 2.678033e-013, 3.285154e-010, -5.150382e-009,
  3.289711e-011, 2.886982e-013, 1.46228e-010, -2.101282e-009,
  7.596613e-011, 1.083126e-013, 2.664249e-010, -3.512665e-009,
  2.988038e-011, 1.966947e-013, 1.721988e-010, -1.644469e-009,
  6.461839e-011, -3.619825e-013, 3.725326e-010, -2.232637e-009,
  2.720721e-011, 1.740702e-013, 8.787672e-011, -1.292279e-009,
  5.529543e-011, -1.726669e-013, 3.173075e-010, -1.173191e-009,
  2.485449e-011, 1.856337e-013, -6.94222e-011, -1.0454e-009,
  4.762206e-011, 9.53694e-014, 1.679692e-010, -4.571889e-010,
  2.277519e-011, 1.861742e-013, 9.091328e-011, -6.845257e-010,
  4.114636e-011, 1.683459e-013, 1.351775e-010, 1.429314e-010,
  2.089262e-011, 1.675215e-013, 3.282472e-011, -3.877256e-010,
  3.562586e-011, 4.262933e-014, 1.003748e-010, 5.042689e-010,
  1.919804e-011, 1.382077e-013, 2.251453e-011, -2.54149e-010,
  3.10947e-011, 1.495005e-014, 1.067664e-010, 8.426829e-010,
  1.764062e-011, 1.361519e-013, -1.097211e-010, -1.768488e-010,
  2.72379e-011, 9.414525e-014, 2.039044e-010, 1.226816e-009,
  1.628732e-011, 1.31162e-013, 9.760202e-011, 1.299755e-010,
  2.386601e-011, 1.684137e-013, -1.476903e-011, 1.284713e-009,
  1.502722e-011, 1.370578e-013, -1.079247e-010, 1.44003e-010,
  2.101066e-011, 1.178166e-013, 1.343749e-010, 1.53653e-009,
  1.389803e-011, 1.208059e-013, -1.433468e-010, 2.163721e-010,
  1.854613e-011, 4.438315e-014, 2.420566e-013, 1.499312e-009,
  1.287296e-011, 1.002387e-013, 7.576488e-012, 3.823121e-010,
  1.63882e-011, -2.180152e-014, -4.261479e-011, 1.548845e-009,
  1.19134e-011, 7.959819e-014, 4.82184e-011, 4.800542e-010,
  1.451339e-011, -7.60117e-014, 1.346128e-010, 1.676413e-009,
  1.104724e-011, 7.029657e-014, 1.012019e-010, 5.977751e-010,
  1.287736e-011, -1.316721e-015, 1.446039e-011, 1.684692e-009,
  1.024938e-011, 9.613409e-014, -1.14711e-010, 5.373039e-010,
  1.144194e-011, 2.123506e-013, 1.64141e-011, 1.704075e-009,
  9.51079e-012, 1.497431e-013, -1.011216e-010, 6.141272e-010,
  1.016868e-011, 2.951804e-013, -1.437801e-010, 1.59815e-009,
  8.824596e-012, 1.690799e-013, 5.036543e-011, 7.490095e-010,
  9.051452e-012, 2.682772e-013, -1.721672e-010, 1.555411e-009,
  8.187271e-012, 1.601054e-013, -8.503767e-011, 7.026859e-010,
  8.06858e-012, 1.19213e-013, 2.208956e-011, 1.618905e-009,
  7.600819e-012, 1.013653e-013, -2.236327e-011, 7.2901e-010,
  7.196191e-012, -1.476994e-013, 1.187338e-011, 1.484425e-009,
  7.061281e-012, 1.107772e-014, 8.647482e-011, 7.888411e-010,
  6.425172e-012, -3.158399e-013, 8.484769e-011, 1.417788e-009,
  6.556616e-012, -4.538347e-014, 1.765615e-010, 8.306844e-010,
  5.745364e-012, -3.181537e-013, 1.265501e-011, 1.3138e-009,
  6.096122e-012, -5.059097e-014, 2.579226e-011, 7.954639e-010,
  5.137946e-012, -2.079934e-013, 7.673933e-011, 1.306429e-009,
  5.676867e-012, -1.17936e-014, 7.924337e-012, 7.411963e-010,
  4.615329e-012, -9.695066e-014, 6.668247e-011, 1.342868e-009,
  5.293036e-012, 3.18464e-014, -5.569571e-011, 6.717936e-010,
  4.137328e-012, -2.597718e-014, 1.761231e-010, 1.382072e-009,
  4.937809e-012, 5.744665e-014, -8.980129e-011, 6.816344e-010,
  3.716155e-012, 2.961723e-015, 8.824103e-011, 1.294919e-009,
  4.609009e-012, 6.736658e-014, -3.377235e-011, 7.515858e-010,
  3.334245e-012, -3.201928e-014, 2.479032e-011, 1.184607e-009,
  4.29603e-012, 4.208465e-014, 3.415802e-011, 7.496462e-010,
  2.980364e-012, -9.406987e-014, -5.20501e-011, 1.054001e-009,
  4.06197e-012, -7.55802e-015, 5.857643e-011, 7.720528e-010,
  2.701874e-012, -1.903456e-013, 6.547055e-011, 1.056132e-009,
  3.761189e-012, -5.717462e-014, -2.07125e-011, 6.519021e-010,
  2.432572e-012, -2.427999e-013, 2.931945e-011, 9.729273e-010,
  3.504873e-012, -8.284223e-014, 1.091847e-010, 7.516331e-010,
  2.198439e-012, -2.601742e-013, 7.853954e-011, 9.748723e-010,
  3.274399e-012, -1.027392e-013, 9.662831e-011, 7.055397e-010,
  1.946211e-012, -2.789156e-013, 1.449718e-010, 9.448567e-010,
  3.087361e-012, -1.310755e-013, 1.877076e-010, 7.655494e-010,
  1.764279e-012, -2.933849e-013, 1.988398e-010, 9.108386e-010,
  2.877626e-012, -1.459811e-013, -7.162008e-012, 6.074524e-010,
  1.618573e-012, -2.898925e-013, 2.59595e-010, 8.861234e-010,
  2.682184e-012, -1.469332e-013, 1.563643e-010, 6.764033e-010,
  1.4637e-012, -2.647472e-013, 1.601958e-010, 8.892874e-010,
  2.512169e-012, -1.339257e-013, 3.08797e-011, 6.464271e-010,
  1.325921e-012, -2.227707e-013, 2.453467e-010, 8.521466e-010,
  2.356376e-012, -1.067364e-013, 4.794168e-011, 6.207563e-010,
  1.198628e-012, -1.433463e-013, 1.233969e-010, 7.686993e-010,
  2.213231e-012, -5.914168e-014, 4.543759e-011, 6.258801e-010,
  1.091131e-012, -9.20184e-014, 7.444635e-011, 7.627776e-010,
  2.080088e-012, -2.82979e-014, 1.004472e-010, 6.714192e-010,
  9.940732e-013, -8.46348e-014, -1.189882e-010, 5.492345e-010,
  1.950848e-012, -2.630735e-014, -7.64581e-011, 5.188868e-010,
  9.014293e-013, -1.302041e-013, 1.009007e-010, 6.276505e-010,
  1.823378e-012, -6.794e-014, 2.55123e-011, 5.433941e-010,
  8.22539e-013, -1.750409e-013, 1.395088e-010, 6.651769e-010,
  1.700729e-012, -1.132493e-013, 1.234947e-010, 6.174707e-010,
  7.439185e-013, -2.304332e-013, 2.03806e-010, 5.888425e-010,
  1.600903e-012, -1.658538e-013, 2.662437e-010, 6.721595e-010,
  6.775736e-013, -2.640723e-013, 4.864509e-011, 4.799655e-010,
  1.499157e-012, -2.054239e-013, 2.867359e-010, 6.203837e-010,
  6.084452e-013, -2.729661e-013, 3.063929e-010, 5.930081e-010,
  1.409567e-012, -2.216733e-013, 1.955057e-010, 5.562495e-010,
  6.076412e-013, -2.946867e-013, 1.385304e-010, 4.256054e-010,
  1.36649e-012, -2.549608e-013, 2.820198e-010, 5.736221e-010,
  5.090655e-013, -2.9893e-013, 2.359266e-010, 4.840432e-010,
  1.243163e-012, -2.683242e-013, 2.90312e-010, 5.278418e-010,
  4.541468e-013, -2.767729e-013, 1.782969e-010, 4.18219e-010,
  1.166731e-012, -2.573217e-013, 3.01819e-010, 5.149493e-010,
  4.158173e-013, -2.15209e-013, 1.456839e-010, 4.248542e-010,
  1.096922e-012, -1.958843e-013, 1.554994e-010, 4.841191e-010,
  3.939366e-013, -1.585819e-013, 1.397673e-010, 4.5103e-010,
  1.092713e-012, -1.515619e-013, -1.001573e-011, 3.711305e-010,
  3.547788e-013, -1.255723e-013, 1.1861e-010, 4.471022e-010,
  9.937263e-013, -1.212389e-013, 9.645993e-011, 4.417108e-010,
  3.182841e-013, -1.213217e-013, 5.409353e-011, 3.653217e-010,
  9.119549e-013, -1.157517e-013, 1.64051e-010, 5.274215e-010,
  2.919132e-013, -1.172936e-013, 1.326594e-010, 3.872055e-010,
  8.59158e-013, -1.140361e-013, 1.722238e-010, 4.645037e-010,
  2.685807e-013, -1.028291e-013, 1.167589e-010, 3.783274e-010,
  8.059365e-013, -1.032599e-013, 6.500376e-011, 3.841661e-010,
  2.455608e-013, -9.665626e-014, 1.685711e-010, 3.889015e-010,
  7.543003e-013, -9.784919e-014, -7.654924e-012, 3.036839e-010,
  2.229456e-013, -9.707607e-014, 2.000945e-010, 3.725495e-010,
  7.075848e-013, -1.057306e-013, 1.216958e-010, 3.933375e-010,
  2.022262e-013, -9.489463e-014, 3.998285e-011, 2.706855e-010,
  6.686734e-013, -1.115054e-013, 2.45448e-010, 4.215418e-010,
  1.850212e-013, -8.069542e-014, 1.051793e-011, 2.256406e-010,
  6.243873e-013, -9.664262e-014, -1.339578e-011, 3.019021e-010,
  1.686799e-013, -6.237892e-014, 1.052296e-010, 3.396725e-010,
  5.846234e-013, -7.465799e-014, 5.851801e-011, 3.62666e-010,
  1.58234e-013, -5.230751e-014, 1.160609e-010, 3.016056e-010,
  5.5458e-013, -6.356006e-014, 5.013805e-011, 3.413234e-010,
  1.485115e-013, -4.232229e-014, 2.37967e-010, 3.944589e-010,
  5.218756e-013, -5.515016e-014, 1.881677e-010, 4.155159e-010,
  1.390158e-013, -4.538444e-014, 5.662286e-011, 2.033141e-010,
  4.920465e-013, -4.436603e-014, 1.237495e-010, 3.355174e-010,
  1.868627e-013, -5.681247e-014, 1.035387e-010, 3.033067e-010,
  4.352551e-013, -4.893652e-014, -1.705698e-011, 2.447422e-010,
  1.20632e-013, -4.602112e-014, 8.249876e-011, 2.464938e-010,
  4.391998e-013, -5.634738e-014, 1.595988e-011, 2.523608e-010,
  1.105992e-013, -4.048434e-014, 4.000061e-011, 2.17523e-010,
  4.149316e-013, -6.645725e-014, 2.131271e-010, 4.108791e-010,
  9.977935e-014, -5.426722e-014, 9.497579e-011, 2.215168e-010,
  3.892539e-013, -8.241712e-014, 1.138102e-010, 3.677384e-010,
  1.61698e-013, -7.408157e-014, 1.015835e-010, 2.082608e-010,
  3.763504e-013, -1.02434e-013, 2.094631e-010, 3.097117e-010,
  1.061125e-013, -7.152761e-014, 8.775923e-011, 2.704078e-010,
  3.48107e-013, -1.125291e-013, 1.318515e-011, 2.417878e-010,
  8.923463e-014, -7.17982e-014, 2.11808e-010, 2.797002e-010,
  3.293483e-013, -1.19342e-013, 3.037193e-011, 1.404994e-010,
  8.195258e-014, -7.194199e-014, 5.780388e-011, 1.013844e-010,
  3.092889e-013, -1.199923e-013, 1.597488e-010, 2.808916e-010,
  7.640671e-014, -6.586057e-014, 5.533341e-011, 1.345277e-010,
  2.927938e-013, -1.194914e-013, 1.438012e-010, 2.531561e-010,
  6.978778e-014, -5.154968e-014, -2.29474e-012, 9.2088e-011,
  2.832328e-013, -9.992841e-014, 1.747288e-010, 2.417508e-010,
  7.514523e-014, -4.236916e-014, -4.849478e-011, 4.876367e-011,
  2.673768e-013, -7.094032e-014, 7.227435e-011, 2.268741e-010,
  7.147624e-014, -2.616592e-014, -1.71463e-011, 4.818044e-011,
  2.470781e-013, -6.937464e-014, 1.117928e-010, 2.02447e-010,
  5.847508e-014, -2.396116e-014, 1.193412e-010, 1.427816e-010,
  2.055302e-013, -5.67724e-014, 2.313219e-011, 1.739626e-010,
  4.621778e-014, -2.53002e-014, 2.297913e-010, 2.871489e-010,
  1.735729e-013, -4.928785e-014, 1.006445e-010, 1.562224e-010,
  5.920187e-014, -2.996249e-014, 4.260679e-011, 1.698458e-010,
  2.138126e-013, -6.006836e-014, 1.362221e-010, 2.860921e-010,
  5.449787e-014, -3.262089e-014, -7.684041e-011, 4.513374e-011,
  1.995148e-013, -6.749196e-014, 6.936296e-011, 1.588022e-010,
  5.494023e-014, -3.495652e-014, -1.034587e-010, 1.040744e-011,
  1.882316e-013, -7.453511e-014, 8.807696e-011, 2.250534e-010,
  6.006143e-014, -3.494121e-014, 7.47209e-011, 1.308559e-010,
  2.506573e-013, -8.573343e-014, 6.404936e-011, 1.730709e-010,
  5.084629e-014, -2.949922e-014, 7.097438e-011, 1.506538e-010,
  1.662735e-013, -6.528874e-014, 1.637885e-010, 2.415165e-010,
  4.988865e-014, -2.377428e-014, 1.057273e-010, 1.407331e-010,
  1.608012e-013, -5.534958e-014, 7.462267e-011, 2.087562e-010,
  4.72714e-014, -2.365876e-014, 2.588733e-011, 9.429574e-011,
  1.519773e-013, -5.56682e-014, 1.023103e-010, 1.683323e-010,
  4.851357e-014, -2.794954e-014, 2.928741e-011, 1.058716e-010,
  1.454112e-013, -6.165465e-014, -1.676222e-012, 8.049391e-011,
  4.553349e-014, -3.088325e-014, 8.231683e-011, 1.387342e-010,
  1.373683e-013, -6.277789e-014, 9.07967e-011, 1.471757e-010,
  4.453908e-014, -2.87735e-014, -7.294125e-011, 3.951283e-011,
  1.277311e-013, -7.066019e-014, 1.361974e-010, 2.068944e-010,
  5.124104e-014, -3.231996e-014, 5.412501e-011, 8.933279e-011,
  1.223568e-013, -7.201728e-014, 7.150708e-012, 1.004375e-010,
  9.2627e-014, -3.54207e-014, 1.507855e-010, 1.59952e-010,
  1.001041e-013, -6.487878e-014, 8.768258e-011, 1.90682e-010,
  6.894772e-014, -2.713025e-014, 6.070502e-011, 1.184546e-010,
  1.036436e-013, -5.551861e-014, 1.011677e-010, 1.475494e-010,
  1.80395e-014, -1.533443e-014, 7.553715e-011, 1.155378e-010,
  5.987168e-014, -4.304776e-014, 1.211731e-010, 2.01827e-010,
  3.785198e-014, -1.564221e-014, 5.850369e-011, 1.341772e-010,
  9.452731e-014, -4.51782e-014, 6.684891e-011, 1.410146e-010,
  7.012705e-014, -2.45181e-014, 7.28254e-011, 1.314921e-010,
  1.030012e-013, -4.613369e-014, 8.011192e-011, 1.317594e-010,
  9.696168e-014, -2.82791e-014, 6.065841e-011, 1.202819e-010,
  1.026177e-013, -4.2625e-014, 4.785723e-011, 1.583282e-010,
  4.425477e-014, -1.925133e-014, 6.954051e-011, 1.504187e-010,
  9.062168e-014, -4.265582e-014, 2.851148e-011, 8.014418e-011,
  4.017366e-014, -2.205779e-014, 1.700103e-010, 1.774839e-010,
  8.246051e-014, -4.301338e-014, 6.306112e-011, 1.860091e-010,
  4.034625e-014, -1.678456e-014, -1.573431e-012, 2.468247e-011,
  8.287234e-014, -3.649142e-014, 1.761184e-010, 2.215281e-010,
  4.125863e-014, -1.254216e-014, 6.93199e-011, 1.196604e-010,
  7.794088e-014, -3.332751e-014, -9.124129e-012, 1.057632e-010,
  3.878809e-014, -1.24099e-014, -3.562109e-011, 1.288824e-011,
  7.578041e-014, -2.871881e-014, -8.282551e-011, 1.387499e-011,
  4.242679e-014, -1.171774e-014, 1.040736e-010, 1.545101e-010,
  6.85378e-014, -2.403193e-014, -9.557196e-011, -4.958707e-012,
  3.602945e-014, -7.417674e-015, -9.8167e-011, -2.711468e-011,
  6.449694e-014, -1.669895e-014, -1.218579e-011, 9.837159e-011,
  2.857588e-014, -2.669116e-015, 5.034151e-011, 1.348466e-010,
  -3.878985e-015, -3.880642e-015, -1.909794e-012, 9.646329e-011,
  4.036513e-014, -8.080818e-015, 3.782307e-011, 8.137598e-011,
  6.564409e-014, -2.127115e-014, 2.942516e-011, 1.126989e-010,
  4.097549e-014, -1.482556e-014, 1.149981e-012, 9.858499e-011,
  5.720844e-014, -2.013972e-014, -1.595452e-011, 9.081743e-011,
  3.747706e-014, -1.388573e-014, -1.567287e-012, 7.511334e-011,
  5.805486e-014, -2.602663e-014, 3.490052e-011, 1.055952e-010,
  2.990876e-014, -1.392481e-014, -1.444516e-010, -1.425264e-010,
  1.143717e-013, -3.869738e-014, 7.497782e-011, 1.181037e-010,
  3.781927e-014, -1.667014e-014, 6.049701e-012, 5.038634e-011,
  7.695641e-014, -3.897052e-014, 4.839057e-011, 1.224028e-010,
  3.750967e-014, -1.89133e-014, 4.705685e-011, -1.372203e-011,
  5.792154e-014, -3.303563e-014, 1.403086e-010, 1.505715e-010,
  3.713163e-014, -1.592359e-014, -3.800404e-011, -4.696809e-011,
  4.232074e-014, -2.334225e-014, 1.985321e-013, 3.501585e-011,
  3.492534e-014, -1.456869e-014, 1.783886e-010, 1.28029e-010,
  4.478556e-014, -2.221463e-014, 2.109886e-010, 1.926475e-010,
  3.750744e-014, -1.139596e-014, 5.158436e-011, 5.249666e-011,
  4.270887e-014, -2.389825e-014, 4.565526e-011, 1.150043e-010,
  3.817552e-014, -1.333323e-014, 5.523309e-012, 7.21289e-011,
  3.90866e-014, -1.75357e-014, -6.838267e-011, 5.339253e-012,
  3.081558e-014, -1.75467e-014, 4.628253e-011, 3.33037e-011,
  3.642737e-014, -1.563514e-014, 3.456476e-011, 4.821146e-011,
  3.878858e-014, -1.522318e-014, -4.513939e-011, -2.897997e-011,
  3.727265e-014, -2.040423e-014, 8.117113e-011, 1.661595e-010,
  9.382875e-014, -2.570148e-014, -1.719264e-011, 2.374446e-011,
  1.640379e-014, -1.624246e-014, -5.307014e-011, 2.349205e-011,
  2.900126e-014, -1.629101e-014, 1.310692e-011, 2.171976e-011,
  3.301868e-014, -2.059287e-014, -5.825229e-011, 9.616705e-012,
  3.192153e-014, -1.684107e-014, 3.045422e-011, 7.043125e-012,
  3.653857e-014, -2.134435e-014, 2.70563e-010, 2.62266e-010,
  3.205369e-014, -1.869887e-014, 1.315911e-010, 8.281565e-011,
  3.450264e-014, -2.296957e-014, 6.699473e-011, 6.677831e-011,
  1.043576e-013, -3.032409e-014, 1.412543e-010, 9.762127e-011,
  5.332376e-014, -2.458907e-014, 1.567135e-010, 1.41479e-010,
  3.353722e-014, -1.476237e-014, 4.571436e-011, 7.493459e-011,
  3.09987e-014, -1.733048e-014, 2.98032e-011, 6.961021e-011,
  2.556485e-014, -1.647183e-014, 5.215471e-011, 3.802421e-011,
  2.709908e-014, -1.267708e-014, 6.983126e-011, 9.812093e-011,
  2.925019e-014, -1.669218e-014, 1.42798e-013, -2.053799e-011,
  2.897086e-014, -1.773274e-014, 9.485018e-012, 6.996528e-011,
  3.137394e-014, -1.631632e-014, 9.515405e-012, 6.222679e-011,
  2.286185e-014, -1.680007e-014, -1.376079e-010, -9.919463e-011,
  3.090567e-014, -1.661278e-014, -5.132328e-011, -6.30245e-012,
  2.285066e-014, -1.258115e-014, 9.223571e-011, 1.083119e-010,
  3.044688e-014, -1.360367e-014, -1.828591e-010, -5.660889e-011,
  2.689601e-014, -1.173091e-014, -4.159544e-011, 1.752694e-011,
  3.304372e-014, -1.342444e-014, -6.558275e-011, 1.329886e-011,
  2.716381e-014, -7.042972e-015, -6.192141e-012, 6.159043e-011,
  3.076701e-014, -7.382152e-015, -4.639916e-011, -3.771331e-012,
  2.544105e-014, -5.234573e-015, -1.622179e-011, 8.458587e-011,
  3.790254e-014, -2.037037e-014, 9.782769e-011, 5.795691e-011,
  2.364116e-014, -1.046363e-014, -8.252414e-011, -5.589307e-011,
  3.411154e-014, -1.249038e-014, -2.151423e-011, 1.388748e-011,
  2.691396e-014, -9.869615e-015, 1.222805e-012, 6.016555e-011,
  2.75837e-014, -6.925163e-015, 5.242612e-011, 9.478776e-011,
  2.769843e-014, -1.978967e-014, -5.479607e-011, -9.02016e-012,
  2.989552e-014, -1.150256e-014, -3.178129e-011, 2.117356e-011,
  3.733928e-015, -8.079676e-015, -1.101325e-011, 3.936092e-011,
  2.238647e-014, -1.37282e-014, -2.244114e-011, -3.518469e-011,
  -3.551461e-014, -2.734966e-015, 1.093602e-011, -9.994824e-012,
  2.52563e-014, -1.228697e-014, -1.712096e-011, 2.726921e-011,
  2.149804e-014, -1.098059e-014, -3.906435e-011, -7.963213e-012,
  2.785589e-014, -1.233084e-014, -6.175688e-011, -1.280467e-011,
  2.261431e-014, -4.199553e-015, 1.910016e-011, 8.153457e-011,
  3.225056e-014, -1.495542e-014, -5.466881e-011, -1.035359e-011,
  1.806406e-014, -5.540692e-015, 1.194027e-010, 1.173318e-010,
  6.746176e-014, -1.82306e-014, 8.95588e-011, 8.141955e-011,
  -4.324944e-014, 3.380249e-015, -8.206629e-011, -1.476329e-011,
  2.600696e-014, -1.113015e-014, 1.839184e-010, 1.579236e-010,
  2.000181e-014, -9.53377e-015, 1.462959e-010, 1.646661e-010,
  2.487317e-014, -1.198896e-014, 3.124652e-011, 3.147125e-011,
  1.980299e-014, -1.241941e-014, 4.125293e-011, 4.939458e-011,
  2.602789e-014, -1.486514e-014, 1.204773e-010, 6.743213e-011,
  2.003191e-014, -1.073521e-014, 1.03871e-010, 3.592537e-011,
  3.133851e-014, -9.533147e-015, -9.246483e-011, -4.888588e-011,
  1.999648e-014, -8.089021e-015, 5.092559e-011, 6.613879e-011,
  2.745176e-014, -4.98064e-015, 5.931305e-012, 6.011978e-011,
  1.502847e-014, -1.844039e-015, 1.468802e-010, 1.228079e-010,
  2.533463e-014, -7.074639e-015, -6.260232e-013, -1.379057e-011,
  1.444467e-014, -5.673802e-015, 5.756651e-012, 7.756885e-011,
  2.756962e-014, -1.1739e-014, 7.771646e-011, 8.964787e-011,
  1.820908e-014, -5.911568e-015, 3.046184e-012, 1.039847e-011,
  -2.583717e-014, -1.992008e-015, -2.007405e-011, 3.134828e-011,
  6.360032e-015, -5.273077e-015, 1.382526e-010, 1.310329e-010,
  1.341235e-014, -8.280632e-015, 5.799158e-012, 3.21266e-011,
  1.33114e-014, -8.81483e-015, 9.945626e-012, 5.900325e-011,
  2.962223e-014, -1.84097e-015, 1.971944e-010, 1.193409e-010,
  1.652064e-014, -7.69184e-015, 1.078187e-010, 1.34401e-010,
  2.979738e-014, -1.037519e-014, 2.605244e-010, 1.217847e-010,
  1.939019e-014, -5.886547e-015, -6.736762e-011, 6.270835e-011,
  5.405537e-014, -1.810353e-014, 2.432154e-011, 7.520862e-012,
  2.586037e-014, -9.598698e-015, 1.954313e-010, 2.048674e-010,
  6.910821e-014, -1.776912e-014, 1.096082e-011, 1.123908e-011,
  3.298427e-014, -1.722948e-014, 7.454908e-011, 9.018354e-012,
  2.001366e-014, -9.697785e-015, 1.153267e-010, 3.728238e-011,
  1.25219e-014, -8.755302e-015, 1.937456e-010, 1.794242e-010,
  1.883868e-014, -1.092744e-014, -1.806254e-010, -1.863001e-010,
  1.502617e-014, -1.099229e-014, 1.904601e-010, 1.330639e-010,
  2.241052e-014, -8.817402e-015, 4.843742e-012, 7.482948e-012,
  7.046077e-015, -1.050813e-014, 3.088832e-012, 4.446145e-011,
  3.052352e-014, -1.338835e-014, -5.949246e-011, 3.912316e-011,
  1.018653e-014, -6.346424e-015, -3.691653e-011, -7.50252e-011,
  2.593432e-014, -1.144389e-014, -1.058886e-011, -1.070018e-011,
  1.240878e-014, -1.531455e-015, -4.719018e-011, -6.640433e-011,
  2.058188e-014, -9.478461e-015, -1.738135e-010, -1.158322e-010,
  1.833261e-014, -6.875662e-015, 5.903774e-011, 6.869703e-011,
  2.692447e-014, -1.450211e-014, -6.308986e-011, -8.80705e-011,
  8.531297e-015, -7.677976e-015, 5.020281e-011, 2.495989e-011,
  2.423478e-014, -1.430656e-014, -9.989613e-011, -8.843219e-011,
  -5.969807e-014, -7.675795e-016, 8.245783e-011, 6.649601e-011,
  2.020286e-014, -1.113209e-014, 6.411304e-011, 8.620426e-011,
  1.341663e-014, -7.663254e-015, 6.569119e-011, 4.760208e-011,
  2.532809e-014, -1.518092e-014, 9.60844e-011, 1.174557e-010,
  6.240964e-015, -6.410642e-015, 6.858571e-012, -6.705154e-012,
  1.975701e-014, -1.190753e-014, 1.00001e-010, 7.757436e-011,
  1.097257e-014, -6.955658e-015, 1.747626e-010, 1.285318e-010,
  6.350865e-014, -1.252356e-014, 1.61466e-010, 1.402782e-010,
  -3.456004e-014, -1.866119e-015, -1.962897e-012, 3.985609e-011,
  2.795234e-014, -1.141872e-014, -1.965711e-011, -2.36071e-011,
  -4.963289e-016, -3.175608e-015, 3.545038e-011, 5.123318e-011,
  1.548905e-014, -1.334636e-014, -1.325051e-011, -6.621127e-013,
  5.634508e-015, -3.179333e-015, -5.748839e-011, -7.991382e-012,
  2.489804e-014, -8.708672e-015, 1.529628e-010, 1.241545e-010,
  7.983299e-015, -9.096485e-015, 1.597818e-012, 2.97525e-011,
  1.588222e-014, -9.369188e-015, 4.255242e-012, 1.206696e-011,
  1.358971e-014, -6.804294e-015, -6.708541e-011, -3.334174e-011,
  1.390381e-014, -8.950695e-015, 2.116497e-011, 1.745688e-011,
  2.209798e-014, -8.267845e-015, 2.834825e-011, 1.658595e-011,
  1.852107e-014, -4.599413e-015, -2.69056e-011, 3.50737e-011,
  1.604055e-014, -2.524328e-015, 5.230463e-012, 3.606157e-011,
  1.338372e-014, -1.49806e-014, -1.53728e-010, -1.003472e-010,
  1.20709e-014, -1.575812e-015, 4.650433e-011, 6.976142e-011,
  2.488941e-014, -1.456058e-014, 3.928813e-011, -2.929229e-011,
  9.332117e-015, -4.166137e-015, 7.546619e-011, 1.299524e-010,
  2.908942e-014, -1.581382e-014, -5.073601e-011, -3.906756e-011,
  1.42126e-014, 3.027228e-015, 1.112801e-011, 7.496023e-011,
  1.870996e-014, -1.280878e-014, 2.14372e-010, 9.259573e-011,
  1.442206e-014, -6.501842e-016, 1.078066e-010, 1.417013e-010,
  7.287566e-015, -9.882481e-015, 1.51908e-010, 1.475151e-010,
  1.136565e-014, -5.189723e-015, 7.341047e-011, 1.000235e-010,
  4.949211e-015, -2.538006e-015, -1.532033e-010, -1.503516e-010,
  3.301969e-015, -1.262392e-015, -2.379359e-010, -1.71226e-010,
  4.76459e-014, 3.317294e-015, -1.787575e-012, 3.420502e-012,
  3.330874e-014, 3.547826e-015, -6.500527e-012, 2.905489e-011,
  5.309826e-014, 3.279984e-015, -2.325577e-011, -8.534407e-012,
  3.175919e-014, 1.995299e-015, 4.89508e-012, 3.726094e-011,
  5.10704e-014, 1.857503e-015, -3.21761e-012, 4.724442e-013,
  1.916608e-014, 4.348045e-015, 9.327792e-013, 3.109776e-011,
  7.434748e-014, -4.352382e-016, -2.833491e-013, 8.216088e-012,
  1.876715e-014, 3.731432e-015, -6.042634e-013, 3.933023e-011,
  5.022101e-014, -1.380665e-015, -1.089948e-012, 3.605634e-012,
  3.718287e-014, 3.158717e-015, 2.252396e-012, 3.320786e-011,
  5.119877e-014, 2.855443e-015, 7.468275e-012, 1.48815e-011,
  3.776953e-014, 3.676358e-015, 3.886672e-012, 2.967118e-011,
  6.244458e-014, -1.669031e-016, -3.789089e-012, 1.30106e-013,
  -3.222114e-014, 1.698138e-014, 4.183513e-012, 4.75612e-011,
  5.559009e-014, 2.721996e-015, -2.623527e-012, 3.571524e-012,
  4.089376e-014, 6.344741e-015, -4.480922e-012, 3.608129e-011,
  5.475166e-014, 3.074781e-015, -3.779699e-012, 1.754141e-012,
  4.197213e-014, 8.281349e-015, -6.457959e-012, 3.592153e-011,
  5.438385e-014, -2.674728e-014, -9.379389e-012, -4.210961e-012,
  3.237838e-014, -1.208465e-014, -7.660964e-012, 3.608651e-011,
  1.264312e-013, -2.751502e-015, -9.93131e-012, -3.191659e-012,
  6.630522e-014, -1.638564e-015, -5.501984e-012, 4.072743e-011,
  6.726031e-014, 8.041414e-017, 2.127284e-012, 3.771767e-012,
  4.888519e-014, 7.032987e-015, -1.811191e-012, 4.581334e-011,
  5.264944e-014, 3.547638e-015, -2.714082e-012, -1.727635e-012,
  7.98586e-014, 4.856994e-015, 7.866702e-013, 4.79924e-011,
  6.181311e-014, 2.315019e-015, 2.60818e-012, 7.516101e-013,
  5.202599e-014, 7.203392e-015, -6.583701e-012, 3.498656e-011,
  6.440425e-014, 2.265598e-015, -2.318057e-012, -2.247573e-012,
  5.007024e-014, 7.359207e-015, -6.958043e-012, 4.413774e-011,
  6.883158e-014, 2.160835e-015, 5.842805e-012, 8.498297e-012,
  4.81604e-014, 5.719228e-015, -9.169078e-013, 4.581793e-011,
  7.52561e-014, 2.407823e-015, -5.473895e-012, -4.679973e-012,
  4.885537e-014, 6.456133e-015, -3.505032e-012, 4.49411e-011,
  7.123468e-014, 2.371097e-015, 1.948428e-012, 5.061728e-012,
  5.465138e-014, 9.555527e-015, -4.578079e-012, 5.342117e-011,
  7.316549e-014, 3.641331e-016, 1.497747e-012, -5.285387e-013,
  5.731762e-014, 1.329484e-014, -4.859402e-012, 5.51307e-011,
  7.814746e-014, 6.004709e-015, 2.9389e-012, 5.460553e-012,
  5.736377e-014, 8.84316e-015, -6.471871e-012, 5.451237e-011,
  7.87847e-014, 7.65884e-016, 4.966306e-012, 4.699481e-012,
  5.943957e-014, 8.166641e-015, -6.872071e-012, 4.737756e-011,
  7.988486e-014, -6.315222e-016, -4.821529e-012, -1.67088e-012,
  5.962066e-014, 4.968753e-015, -1.925877e-012, 5.415516e-011,
  8.639304e-014, -3.287814e-015, -3.894145e-012, 3.902244e-013,
  5.234826e-014, 3.775549e-015, -1.480563e-011, 4.581826e-011,
  4.715807e-014, 4.184655e-016, -2.454182e-012, 4.476549e-012,
  -1.368321e-014, 1.25361e-014, -4.73182e-012, 4.932101e-011,
  8.80611e-014, -1.328818e-015, 4.20882e-012, 9.078578e-012,
  6.423461e-014, 5.508879e-015, 6.607536e-012, 6.558075e-011,
  9.289754e-014, -2.193227e-015, -3.976795e-012, 4.44396e-012,
  6.465471e-014, 1.982824e-015, 8.385529e-012, 7.169463e-011,
  9.333524e-014, -1.016378e-014, 6.393055e-012, 1.76572e-011,
  6.712456e-014, 2.066746e-015, 6.352628e-012, 6.887804e-011,
  1.673762e-013, -2.079973e-014, -9.01779e-013, 7.305581e-012,
  1.181105e-013, -5.836345e-015, 9.47478e-014, 6.26463e-011,
  1.022272e-013, -1.193425e-014, 2.062184e-012, 1.016896e-011,
  6.530492e-014, -1.120709e-015, -3.591303e-012, 6.526263e-011,
  1.038969e-013, -1.181023e-014, 1.852234e-011, 1.913408e-011,
  7.061511e-014, -2.760534e-015, 4.619947e-012, 7.276241e-011,
  1.062114e-013, -1.301382e-014, 2.072313e-012, 7.101334e-012,
  7.337335e-014, -3.863333e-015, 5.883998e-012, 7.458327e-011,
  1.092065e-013, -1.278079e-014, -4.680962e-012, 1.4955e-011,
  7.60353e-014, 3.104999e-016, 5.135892e-012, 2.538283e-011,
  1.107635e-013, -1.002374e-014, -1.140374e-011, 2.983839e-012,
  7.657177e-014, -3.817744e-015, 6.079817e-012, 7.6012e-011,
  1.125147e-013, -8.410445e-015, -2.423913e-013, 4.24089e-012,
  8.281241e-014, -1.807504e-015, 2.706993e-012, 7.890889e-011,
  1.217194e-013, -9.509558e-015, -6.354446e-012, 5.749771e-012,
  8.195719e-014, 1.538123e-016, -1.109887e-012, 8.282057e-011,
  1.257797e-013, -1.183571e-014, -3.853886e-012, 4.234156e-012,
  7.589738e-014, 1.972157e-015, -5.204368e-012, 7.657122e-011,
  1.180787e-013, -1.591234e-014, 1.491175e-012, -3.666232e-014,
  6.840621e-014, 2.080475e-015, -5.700708e-012, 8.175111e-011,
  1.367436e-013, -1.706798e-014, 4.31321e-012, 5.609748e-012,
  8.694676e-014, -2.367917e-015, -3.370609e-013, 9.044367e-011,
  1.46076e-013, -1.288408e-014, -3.761489e-012, 3.749493e-012,
  9.739976e-014, 2.48573e-017, -1.135824e-012, 9.531473e-011,
  1.431456e-013, -4.310721e-015, -1.309486e-012, 8.915832e-012,
  1.041541e-013, 3.7535e-015, 2.039011e-012, 1.046576e-010,
  1.531519e-013, -4.639879e-016, -4.596083e-012, 5.253981e-012,
  1.461761e-013, -1.797375e-015, 2.119076e-013, 1.12361e-010,
  1.510666e-013, 7.205631e-017, 1.714797e-012, 6.59967e-012,
  9.412504e-014, 9.718911e-015, -5.102363e-012, 1.112937e-010,
  1.562382e-013, 2.265903e-015, -4.32825e-012, -4.891324e-014,
  9.987197e-014, 1.26695e-014, -8.770169e-012, 1.134417e-010,
  1.592544e-013, 4.764296e-015, 3.501278e-012, 1.116033e-011,
  1.003671e-013, 1.388724e-014, -1.057728e-011, 1.184067e-010,
  8.698285e-014, 1.945207e-014, -1.683135e-012, 4.58783e-012,
  9.230188e-014, 1.782173e-014, -7.965639e-012, 1.26669e-010,
  1.712297e-013, 1.17648e-014, -2.40131e-013, 3.974932e-012,
  1.030428e-013, 2.136448e-014, -1.264191e-011, 1.288953e-010,
  1.790745e-013, 1.586116e-014, 1.718268e-012, 1.258347e-011,
  1.065363e-013, 2.037844e-014, -1.399114e-011, 1.360201e-010,
  1.825006e-013, 1.931043e-014, -3.805179e-012, 9.624778e-012,
  1.103294e-013, 2.433852e-014, -2.358785e-011, 1.319339e-010,
  2.0537e-013, 2.148221e-014, 8.204494e-012, 2.744441e-011,
  1.273914e-013, 5.422266e-014, -2.588654e-011, 1.419538e-010,
  1.959895e-013, 3.452257e-014, 6.957354e-012, 1.576928e-011,
  1.131338e-013, 3.248634e-014, -2.98839e-011, 1.475501e-010,
  1.989957e-013, 3.454873e-014, -8.096344e-012, 2.940734e-012,
  1.159899e-013, 3.446583e-014, -3.295377e-011, 1.527239e-010,
  2.045181e-013, 2.74566e-014, 3.703896e-012, 1.96427e-011,
  1.170677e-013, 3.237621e-014, -2.46939e-011, 1.660388e-010,
  2.501474e-013, 1.568082e-014, 1.613249e-012, 1.883529e-011,
  1.069119e-013, 3.157319e-014, -3.260195e-011, 1.636398e-010,
  2.487548e-013, 1.563217e-014, -5.150404e-012, 9.257626e-012,
  1.121649e-013, 2.969683e-014, -3.077504e-011, 1.737161e-010,
  2.306548e-013, 1.718874e-014, 4.644406e-012, 2.223482e-011,
  1.284364e-013, 2.436858e-014, -2.078345e-011, 1.853733e-010,
  2.362105e-013, 1.060854e-014, -1.40453e-013, 1.97287e-011,
  1.309161e-013, 2.125016e-014, -1.657334e-011, 1.916069e-010,
  2.490535e-013, 5.97285e-015, -4.065068e-013, 2.338232e-011,
  1.56206e-013, 1.631247e-014, -1.480001e-011, 2.028081e-010,
  2.679338e-013, 5.71727e-015, -9.022207e-012, 1.892381e-011,
  1.90469e-013, 7.978581e-015, 2.68363e-012, 2.325775e-010,
  2.582076e-013, -8.584461e-016, -1.662654e-012, 3.257208e-011,
  1.390886e-013, 1.372265e-014, -1.593872e-012, 2.320309e-010,
  2.655012e-013, -6.26372e-015, 3.227603e-012, 3.335135e-011,
  1.450418e-013, 1.071985e-014, -3.093717e-012, 2.382108e-010,
  2.714427e-013, -1.362971e-014, 1.376847e-012, 3.369711e-011,
  1.495851e-013, 9.340309e-015, 3.429162e-012, 2.4909e-010,
  2.764756e-013, -1.799021e-014, -4.053814e-013, 3.743934e-011,
  1.527524e-013, 5.649133e-015, 7.662807e-012, 2.623402e-010,
  2.851146e-013, -1.979697e-014, -1.743029e-012, 3.886549e-011,
  1.572804e-013, 5.207405e-015, 9.809047e-012, 2.789905e-010,
  2.925881e-013, -1.7168e-014, 1.561078e-012, 5.080524e-011,
  1.626805e-013, 3.68406e-015, 6.651351e-012, 2.92998e-010,
  2.986928e-013, -1.790847e-014, 1.587561e-012, 5.474477e-011,
  1.704144e-013, 5.673566e-015, 1.65212e-012, 3.03272e-010,
  2.805715e-013, -1.903243e-014, 6.741936e-012, 6.243635e-011,
  1.786045e-013, 3.74535e-015, 5.771553e-012, 3.262912e-010,
  3.084918e-013, -2.542549e-014, 5.582261e-012, 6.216755e-011,
  1.857907e-013, 5.091274e-015, 1.149439e-011, 3.369159e-010,
  3.132186e-013, -2.379824e-014, 7.968692e-012, 7.469759e-011,
  1.942534e-013, 7.333399e-015, 7.026808e-012, 3.513785e-010,
  3.175826e-013, -2.122373e-014, 2.750984e-011, 1.091051e-010,
  2.005108e-013, 1.273519e-014, 3.963768e-012, 3.71151e-010,
  3.818877e-013, -2.398228e-014, 1.138427e-011, 9.910548e-011,
  2.153856e-013, 1.745475e-014, 5.125114e-012, 3.965761e-010,
  3.432919e-013, -1.826237e-014, 1.226957e-011, 1.106162e-010,
  2.277276e-013, 1.480257e-014, 2.11926e-012, 4.125338e-010,
  3.306446e-013, -1.762057e-014, 5.134757e-012, 1.145045e-010,
  2.448221e-013, 1.423145e-014, 1.364007e-011, 4.460376e-010,
  3.320602e-013, -1.967171e-014, 1.845536e-012, 1.238737e-010,
  2.636626e-013, 1.00444e-014, 1.768787e-011, 4.689976e-010,
  3.098832e-013, -2.281373e-014, 8.980737e-012, 1.419223e-010,
  2.595421e-013, 1.284317e-014, 1.45584e-011, 4.855548e-010,
  2.946415e-013, -1.403764e-014, 8.618509e-012, 1.581246e-010,
  2.752127e-013, 2.060483e-014, 4.499056e-012, 5.048117e-010,
  3.310976e-013, -1.292298e-014, 7.50648e-012, 1.753212e-010,
  3.345111e-013, 2.560125e-014, -2.402776e-012, 5.331036e-010,
  3.280669e-013, -3.992819e-015, 4.035206e-012, 1.896655e-010,
  3.670506e-013, 3.503625e-014, -3.335716e-012, 5.695358e-010,
  3.222843e-013, -1.08761e-014, 5.983946e-012, 2.140257e-010,
  4.035778e-013, 3.147786e-014, -8.742199e-012, 5.847995e-010,
  3.167828e-013, -2.105309e-014, 4.242176e-012, 2.387479e-010,
  4.465435e-013, 1.60415e-014, 4.984891e-013, 6.105307e-010,
  3.147936e-013, -2.819652e-014, 6.618861e-012, 2.601352e-010,
  4.958454e-013, 6.305427e-015, 2.146772e-011, 6.468353e-010,
  3.083778e-013, -2.543803e-014, 1.752147e-011, 3.012391e-010,
  5.520235e-013, 8.547071e-015, 2.061419e-011, 6.819046e-010,
  3.015385e-013, -1.045901e-014, 5.319758e-012, 3.219318e-010,
  6.214091e-013, 2.476669e-014, 1.448685e-011, 7.181442e-010,
  3.140487e-013, -4.223444e-015, -8.070431e-013, 3.550063e-010,
  6.831692e-013, 4.042053e-014, -1.244002e-011, 7.345651e-010,
  2.870087e-013, -5.636526e-015, 2.653427e-012, 3.950539e-010,
  7.912712e-013, 2.707883e-014, 6.501989e-012, 7.887224e-010,
  2.826347e-013, -1.470157e-014, 1.874107e-011, 4.539648e-010,
  8.968788e-013, 1.372984e-014, 3.225276e-012, 8.064636e-010,
  2.780925e-013, -1.857233e-014, 3.37086e-012, 4.797024e-010,
  1.020387e-012, 7.554979e-017, 1.740937e-011, 8.539404e-010,
  2.228203e-013, -1.37458e-014, 1.05371e-011, 5.415164e-010,
  1.20701e-012, -1.347584e-014, 3.01948e-011, 8.894883e-010,
  2.647003e-013, -1.910563e-014, 1.818698e-011, 6.04181e-010,
  1.342459e-012, -9.348072e-015, 3.782045e-011, 9.262145e-010,
  2.749761e-013, -2.774798e-014, 2.315687e-011, 6.654553e-010,
  1.528645e-012, -2.734142e-014, 3.380667e-011, 9.476352e-010,
  2.837666e-013, -4.656279e-014, 2.227387e-011, 7.303247e-010,
  1.754406e-012, -5.56994e-014, 5.317291e-011, 9.866613e-010,
  2.802252e-013, -5.642235e-014, 2.755297e-011, 7.989326e-010,
  1.971191e-012, -7.476249e-014, 6.931151e-011, 1.015849e-009,
  3.150555e-013, -4.195908e-014, 3.314133e-011, 8.905575e-010,
  2.289405e-012, -6.220577e-014, 5.338397e-011, 1.043712e-009,
  3.753563e-013, -2.117596e-014, 1.210686e-011, 9.635215e-010,
  2.65987e-012, -3.791221e-014, 2.986191e-011, 1.057224e-009,
  4.398714e-013, -5.218265e-015, 1.331724e-011, 1.063205e-009,
  3.062012e-012, -2.804967e-014, 1.324944e-011, 1.073607e-009,
  5.30772e-013, -1.984533e-014, 2.200435e-011, 1.163173e-009,
  3.525561e-012, -5.272613e-014, 2.696737e-011, 1.095665e-009,
  6.619451e-013, -3.936308e-014, 3.158872e-011, 1.270145e-009,
  4.048403e-012, -9.192017e-014, 3.870406e-011, 1.100628e-009,
  8.264724e-013, -4.288009e-014, 3.831851e-011, 1.385126e-009,
  4.654061e-012, -1.014395e-013, 4.396413e-011, 1.098353e-009,
  1.052057e-012, -1.208965e-014, 2.278603e-011, 1.507472e-009,
  5.346833e-012, -7.50454e-014, 2.910447e-011, 1.092878e-009,
  1.342676e-012, 6.179706e-015, 9.660544e-012, 1.62063e-009,
  6.138816e-012, -6.518242e-014, 1.059561e-011, 1.060389e-009,
  1.716261e-012, 9.114343e-015, 1.715496e-011, 1.747345e-009,
  7.053196e-012, -8.273268e-014, 2.233849e-011, 1.026183e-009,
  2.199175e-012, 7.077114e-014, -8.769879e-012, 1.867181e-009,
  8.113457e-012, -3.054512e-014, -1.155225e-011, 9.540243e-010,
  2.811897e-012, 1.370009e-013, -3.181526e-011, 1.995933e-009,
  9.315616e-012, 2.544342e-014, -4.286553e-011, 8.691846e-010,
  3.594493e-012, 1.478808e-013, -3.087607e-011, 2.123823e-009,
  1.070266e-011, 2.244764e-014, -5.089883e-011, 7.526398e-010,
  4.574239e-012, 1.08674e-013, -3.387819e-011, 2.211368e-009,
  1.231971e-011, -2.353652e-014, -3.08721e-011, 6.102305e-010,
  5.805296e-012, 8.908188e-014, -2.037961e-011, 2.313976e-009,
  1.415265e-011, -4.058262e-014, -5.223987e-011, 4.108785e-010,
  7.381369e-012, 6.610282e-014, -6.592077e-012, 2.408192e-009,
  1.633763e-011, -6.024295e-014, -2.299892e-011, 2.081733e-010,
  9.359874e-012, 4.546234e-014, -9.196953e-012, 2.44772e-009,
  1.876041e-011, -6.263557e-014, -2.642224e-011, -1.01877e-010,
  1.184657e-011, -1.351071e-013, 2.695711e-011, 2.459877e-009,
  2.160897e-011, -1.63886e-013, 7.116627e-012, -4.460088e-010,
  1.496635e-011, -4.068956e-013, 7.738077e-011, 2.3709e-009,
  2.490085e-011, -3.174238e-013, 3.947475e-011, -8.876985e-010,
  1.888234e-011, -4.442805e-013, 7.45849e-011, 2.22766e-009,
  2.866292e-011, -3.170342e-013, 4.06149e-011, -1.406396e-009,
  2.384601e-011, -4.961014e-013, 7.340038e-011, 1.956137e-009,
  3.305144e-011, -3.137867e-013, 3.078958e-011, -2.036246e-009,
  3.010397e-011, -7.638262e-013, 1.13657e-010, 1.535257e-009,
  3.808829e-011, -4.045429e-013, 5.132523e-011, -2.777787e-009,
  3.811614e-011, -1.308891e-012, 1.874755e-010, 8.694314e-010,
  4.397386e-011, -5.826704e-013, 9.997571e-011, -3.698067e-009,
  4.827232e-011, -1.8961e-012, 2.50045e-010, -1.128862e-010,
  5.077244e-011, -7.317899e-013, 1.381872e-010, -4.795563e-009,
  6.136348e-011, -2.650183e-012, 3.39187e-010, -1.525875e-009,
  5.881469e-011, -8.77149e-013, 1.801026e-010, -6.138972e-009,
  7.828065e-011, -3.314179e-012, 3.832293e-010, -3.53096e-009,
  6.828405e-011, -9.091177e-013, 2.076583e-010, -7.752443e-009,
  1.004835e-010, -4.97433e-012, 5.57292e-010, -6.302782e-009,
  7.933858e-011, -1.123648e-012, 2.992129e-010, -9.699399e-009,
  1.294714e-010, -7.136925e-012, 7.318026e-010, -1.014062e-008,
  9.235478e-011, -1.355035e-012, 3.904166e-010, -1.203201e-008,
  1.671456e-010, -8.661103e-012, 7.038483e-010, -1.551314e-008,
  1.059573e-010, -1.499471e-012, 3.666014e-010, -1.488536e-008,
  2.216243e-010, -1.067273e-011, 7.642215e-010, -2.312666e-008,
  1.241102e-010, -1.060951e-012, 3.984123e-010, -1.836769e-008,
  2.950881e-010, -1.481362e-011, 1.047968e-009, -3.405364e-008,
  1.47762e-010, -1.231431e-012, 5.555981e-010, -2.268909e-008,
  4.016565e-010, -1.881508e-011, 1.213618e-009, -5.015981e-008,
  1.759163e-010, -9.883494e-013, 6.488551e-010, -2.812487e-008,
  5.580301e-010, -2.319951e-011, 1.301177e-009, -7.400404e-008,
  2.106498e-010, -6.480067e-013, 7.076168e-010, -3.489594e-008,
  8.033185e-010, -2.838985e-011, 1.517357e-009, -1.114376e-007,
  2.556788e-010, 1.714307e-014, 7.885093e-010, -4.371737e-008,
  1.206849e-009, -3.389894e-011, 2.395282e-009, -1.721707e-007,
  3.152706e-010, 1.594848e-012, 1.107407e-009, -5.529536e-008,
  1.915654e-009, -5.331742e-011, 5.829981e-009, -2.809185e-007,
  3.956186e-010, 4.0872e-012, 1.89764e-009, -7.154443e-008,
  3.163995e-009, -1.052631e-010, 1.454405e-008, -4.979696e-007,
  5.048408e-010, 8.087101e-012, 3.424547e-009, -9.544645e-008,
  4.352048e-009, -2.593176e-010, 3.96635e-008, -1.005409e-006,
  5.982417e-010, 1.306731e-011, 6.285362e-009, -1.333436e-007,
  -7.641501e-010, -5.61224e-010, 1.092542e-007, -2.188767e-006,
  5.229455e-010, 1.954486e-011, 1.091543e-008, -1.848843e-007,
  -1.051183e-008, -5.904491e-010, 1.704322e-007, -3.58243e-006,
  5.651913e-010, 2.64811e-011, 1.25079e-008, -2.206573e-007,
  -1.251003e-008, -5.8653e-010, 1.687414e-007, -3.996301e-006,
  6.244956e-010, 1.527587e-011, 1.018439e-008, -2.229892e-007,
  -9.521573e-009, -1.008693e-009, 1.150235e-007, -3.371832e-006,
  7.114277e-010, -6.889417e-012, 6.906258e-009, -1.905669e-007,
  6.64022e-010, -1.086108e-009, 4.931967e-008, -1.946853e-006,
  7.546916e-010, 3.321087e-013, 4.611865e-009, -1.414135e-007,
  4.405495e-009, -4.342789e-010, 1.871376e-008, -8.950659e-007,
  5.793906e-010, 7.641017e-012, 2.991712e-009, -1.082348e-007,
  3.009442e-009, -8.994212e-011, 6.728921e-009, -4.550708e-007,
  4.571636e-010, 4.845075e-012, 1.544836e-009, -8.36323e-008,
  1.818562e-009, -1.546217e-011, 1.996731e-009, -2.629003e-007,
  3.661698e-010, 1.230357e-012, 6.575624e-010, -6.542239e-008,
  1.151443e-009, -2.011747e-011, 1.077966e-009, -1.63738e-007,
  2.961317e-010, -8.393157e-013, 4.65457e-010, -5.179971e-008,
  7.743657e-010, -2.675919e-011, 1.148524e-009, -1.075676e-007,
  2.43574e-010, -2.356016e-012, 5.91262e-010, -4.156301e-008,
  5.444051e-010, -3.059861e-011, 1.709515e-009, -7.304417e-008,
  2.029428e-010, -2.733532e-012, 8.345898e-010, -3.369559e-008,
  3.944516e-010, -2.487942e-011, 1.786575e-009, -5.051217e-008,
  1.70896e-010, -2.390714e-012, 8.666319e-010, -2.748613e-008,
  2.933533e-010, -1.607209e-011, 1.500785e-009, -3.533554e-008,
  1.452189e-010, -1.721088e-012, 7.248429e-010, -2.257039e-008,
  2.22236e-010, -8.955673e-012, 1.107369e-009, -2.469652e-008,
  1.239913e-010, -1.168879e-012, 5.467732e-010, -1.860448e-008,
  1.702856e-010, -7.744579e-012, 1.090312e-009, -1.717433e-008,
  1.062406e-010, -1.364298e-012, 5.614622e-010, -1.529823e-008,
  1.326003e-010, -6.09995e-012, 1.055851e-009, -1.181694e-008,
  9.278156e-011, -1.062493e-012, 5.643302e-010, -1.25805e-008,
  1.037128e-010, -5.451073e-012, 1.023345e-009, -7.927565e-009,
  8.016757e-011, -1.056401e-012, 5.747095e-010, -1.032243e-008,
  8.16562e-011, -3.989947e-012, 8.545986e-010, -5.059918e-009,
  6.938313e-011, -7.62191e-013, 5.185976e-010, -8.383196e-009,
  6.450104e-011, -1.949139e-012, 5.56029e-010, -2.919754e-009,
  6.013999e-011, -2.141402e-013, 3.613488e-010, -6.783826e-009,
  5.114434e-011, -2.866071e-014, 2.374331e-010, -1.351975e-009,
  5.213387e-011, 2.691859e-013, 1.618385e-010, -5.435949e-009,
  4.063482e-011, -8.687835e-014, 2.182458e-010, -1.958199e-010,
  4.525158e-011, 1.235175e-013, 1.612468e-010, -4.30129e-009,
  3.233342e-011, -5.221095e-013, 2.588585e-010, 6.322676e-010,
  3.934584e-011, -5.657e-014, 2.004504e-010, -3.335891e-009,
  2.577366e-011, -3.2689e-013, 1.90931e-010, 1.204628e-009,
  3.428184e-011, 1.674432e-014, 1.63153e-010, -2.539511e-009,
  2.062536e-011, -6.460894e-014, 1.421297e-010, 1.596415e-009,
  2.99509e-011, 1.245688e-013, 8.780816e-011, -1.901987e-009,
  1.647465e-011, 1.591082e-014, 9.229129e-011, 1.824051e-009,
  2.615597e-011, 1.472127e-013, 7.981218e-011, -1.341238e-009,
  1.313376e-011, -6.604649e-014, 8.56729e-011, 1.981014e-009,
  2.291296e-011, 5.443227e-014, 7.970349e-011, -8.923656e-010,
  1.054479e-011, -7.085727e-014, 6.317283e-011, 2.049825e-009,
  2.001162e-011, 4.58435e-014, 5.798752e-011, -5.197341e-010,
  8.462184e-012, 1.528438e-015, 1.927014e-011, 2.054319e-009,
  1.756889e-011, 7.781472e-014, 3.933548e-011, -1.989263e-010,
  6.749435e-012, 7.223407e-014, 1.073693e-011, 2.040351e-009,
  1.538568e-011, 1.109962e-013, 2.412712e-011, 5.611183e-011,
  5.388238e-012, 4.49502e-014, 2.222329e-011, 2.008997e-009,
  1.350589e-011, 7.63354e-014, 2.037757e-011, 2.632367e-010,
  4.298601e-012, 2.542563e-015, 3.024848e-011, 1.943152e-009,
  1.18679e-011, 3.590882e-014, 5.634707e-012, 4.145115e-010,
  3.424666e-012, -3.676783e-014, 4.049173e-011, 1.858606e-009,
  1.041087e-011, -4.436484e-015, 2.671791e-011, 5.623511e-010,
  2.717232e-012, -6.980699e-014, 2.977808e-011, 1.752421e-009,
  9.141329e-012, -3.547423e-014, 2.808837e-011, 6.642513e-010,
  2.147546e-012, -2.891894e-014, 8.411339e-012, 1.654496e-009,
  8.029801e-012, 7.777114e-015, 2.530872e-011, 7.622404e-010,
  1.700092e-012, 8.512482e-014, -3.489803e-011, 1.547317e-009,
  7.051865e-012, 1.305808e-013, -4.459792e-011, 8.173465e-010,
  1.339437e-012, 1.265637e-013, -4.354112e-011, 1.455263e-009,
  6.185193e-012, 1.756107e-013, -7.381255e-011, 8.660771e-010,
  1.060185e-012, 1.115323e-013, -3.321289e-011, 1.365375e-009,
  5.422122e-012, 1.565504e-013, -6.531722e-011, 9.021265e-010,
  8.398651e-013, 4.824371e-014, -2.105445e-011, 1.25959e-009,
  4.758879e-012, 7.274398e-014, -2.168141e-011, 9.248431e-010,
  6.685327e-013, -6.869004e-014, 3.145245e-011, 1.175954e-009,
  4.172009e-012, -7.791602e-014, 6.512295e-011, 9.403841e-010,
  5.37397e-013, -1.34783e-013, 5.093266e-011, 1.082352e-009,
  3.657794e-012, -1.706433e-013, 1.218685e-010, 9.573961e-010,
  4.332387e-013, -1.348089e-013, 7.949272e-011, 1.015208e-009,
  3.208473e-012, -1.707415e-013, 9.164305e-011, 9.190036e-010,
  3.579824e-013, -8.736581e-014, 4.714572e-011, 9.385323e-010,
  2.818204e-012, -1.111184e-013, 7.561933e-011, 9.331734e-010,
  2.777925e-013, -3.676986e-014, 3.279531e-011, 8.616783e-010,
  2.488018e-012, -4.865282e-014, 4.613385e-011, 9.198329e-010,
  2.628114e-013, -1.091657e-014, 1.998036e-011, 7.895492e-010,
  2.17493e-012, -1.420818e-014, 1.527686e-011, 8.909799e-010,
  2.412345e-013, -3.238501e-015, -6.23674e-012, 7.173221e-010,
  1.912277e-012, 1.321689e-016, 2.879307e-011, 8.908322e-010,
  2.272931e-013, -6.390289e-015, 1.516464e-011, 6.704698e-010,
  1.683649e-012, -1.664769e-014, 2.856756e-012, 8.414525e-010,
  2.747476e-013, -3.73286e-014, 1.720521e-011, 6.049784e-010,
  1.453701e-012, -4.372807e-014, 4.219017e-011, 8.377558e-010,
  2.27642e-013, -5.684389e-014, 1.726677e-011, 5.432521e-010,
  1.302676e-012, -9.038199e-014, 6.068948e-011, 8.050745e-010,
  2.164278e-013, -7.035309e-014, 1.589535e-011, 4.906871e-010,
  1.153946e-012, -1.15018e-013, 7.825126e-011, 7.760318e-010,
  2.187309e-013, -7.597553e-014, 2.61697e-011, 4.589064e-010,
  1.022166e-012, -1.20283e-013, 9.256546e-011, 7.509063e-010,
  2.372682e-013, -8.268075e-014, 4.527266e-011, 4.345821e-010,
  9.495568e-013, -1.301815e-013, 9.269684e-011, 7.255606e-010,
  2.397805e-013, -8.722013e-014, 4.48054e-011, 4.001759e-010,
  8.264876e-013, -1.318315e-013, 1.058091e-010, 6.990613e-010,
  2.34551e-013, -8.381064e-014, 4.829514e-011, 3.543725e-010,
  7.067608e-013, -1.239954e-013, 1.039151e-010, 6.623475e-010,
  2.502475e-013, -7.891398e-014, 3.737525e-011, 3.194205e-010,
  6.38163e-013, -1.111693e-013, 7.96145e-011, 6.240818e-010,
  2.543194e-013, -5.921194e-014, 1.711685e-011, 2.897986e-010,
  5.72822e-013, -8.910322e-014, 7.822051e-011, 6.281629e-010,
  2.557083e-013, -3.483374e-014, -1.655411e-011, 2.429397e-010,
  5.082352e-013, -5.577213e-014, 8.157337e-011, 6.429211e-010,
  2.689884e-013, -1.600653e-014, -4.477407e-012, 2.330799e-010,
  4.613293e-013, -3.574162e-014, 4.55067e-011, 5.960195e-010,
  2.765843e-013, -1.737604e-014, -2.506501e-011, 1.916632e-010,
  4.163391e-013, -3.762996e-014, 4.066118e-011, 5.715052e-010,
  2.811086e-013, -3.967824e-014, 1.249237e-011, 2.140828e-010,
  3.758019e-013, -5.36217e-014, 3.857771e-011, 5.215848e-010,
  2.896807e-013, -5.519052e-014, 9.131185e-012, 1.954534e-010,
  3.158953e-013, -6.576343e-014, 5.747341e-011, 5.012522e-010,
  2.816146e-013, -7.479619e-014, 1.258393e-011, 1.621278e-010,
  3.082648e-013, -8.514093e-014, 1.032546e-010, 4.907819e-010,
  2.841269e-013, -9.422474e-014, 1.963026e-011, 1.640129e-010,
  2.860234e-013, -9.820871e-014, 1.034533e-010, 4.454873e-010,
  2.861405e-013, -1.007998e-013, -6.938635e-013, 1.202757e-010,
  2.616505e-013, -1.030424e-013, 8.435939e-011, 4.243169e-010,
  2.504158e-013, -1.092184e-013, 2.196776e-011, 1.293767e-010,
  3.025537e-013, -1.16498e-013, 1.273211e-010, 4.231889e-010,
  2.77329e-013, -1.258545e-013, 1.520869e-011, 1.164803e-010,
  2.276718e-013, -1.122591e-013, 1.320875e-010, 3.965767e-010,
  2.75485e-013, -1.224861e-013, 1.238223e-013, 9.270747e-011,
  2.082534e-013, -1.033928e-013, 1.13746e-010, 3.717378e-010,
  2.775002e-013, -9.31885e-014, 1.978421e-011, 1.028687e-010,
  1.954373e-013, -7.676574e-014, 9.764066e-011, 3.595223e-010,
  2.324393e-013, -6.240379e-014, 8.944593e-012, 9.012376e-011,
  1.5118e-013, -5.192173e-014, 6.738422e-011, 3.382593e-010,
  2.574965e-013, -5.556504e-014, 2.074178e-011, 9.00708e-011,
  1.670962e-013, -4.576797e-014, 7.604942e-011, 3.602612e-010,
  2.673142e-013, -5.646031e-014, -2.753441e-012, 6.875554e-011,
  1.670329e-013, -4.553592e-014, 7.170977e-011, 3.380622e-010,
  2.658262e-013, -5.746464e-014, 1.319777e-011, 7.162737e-011,
  1.57231e-013, -4.35391e-014, 5.502092e-011, 3.027499e-010,
  2.598534e-013, -5.113921e-014, 6.528545e-012, 6.414928e-011,
  1.506165e-013, -3.951269e-014, 5.278379e-011, 2.808434e-010,
  2.575515e-013, -4.578879e-014, -8.267057e-013, 5.62522e-011,
  1.44321e-013, -3.657204e-014, 4.021062e-011, 2.771209e-010,
  2.520257e-013, -5.181345e-014, -3.670614e-012, 4.486442e-011,
  1.354239e-013, -3.757511e-014, 4.111091e-011, 2.55751e-010,
  2.461212e-013, -5.555971e-014, 2.238492e-012, 4.653951e-011,
  1.294838e-013, -4.157975e-014, 4.140539e-011, 2.398467e-010,
  2.428189e-013, -4.610455e-014, 1.30385e-011, 4.863332e-011,
  1.311361e-013, -3.522693e-014, 4.348128e-011, 2.503443e-010,
  2.398453e-013, -3.645907e-014, -4.417476e-012, 2.856936e-011,
  1.495912e-013, -3.164809e-014, 6.58924e-011, 2.64014e-010,
  2.329154e-013, -3.183279e-014, -1.087245e-011, 1.40237e-011,
  1.167976e-013, -2.129357e-014, 3.173704e-011, 2.383079e-010,
  2.289356e-013, -2.529078e-014, -1.340755e-011, 1.790725e-011,
  1.142022e-013, -1.730687e-014, 2.061091e-011, 2.194769e-010,
  2.219595e-013, -2.275999e-014, 1.366404e-011, 2.627698e-011,
  1.134965e-013, -1.570294e-014, 4.003744e-011, 2.195397e-010,
  2.102836e-013, -2.593276e-014, 1.781542e-011, 4.975592e-011,
  4.01984e-014, -1.104778e-014, 2.675328e-011, 2.102669e-010,
  2.120679e-013, -3.294287e-014, 3.624692e-011, 3.282575e-011,
  1.065675e-013, -2.140134e-014, 3.6374e-011, 2.152001e-010,
  2.061364e-013, -4.286219e-014, 9.340279e-012, 3.797683e-011,
  1.058474e-013, -2.543857e-014, 5.60684e-011, 2.007212e-010,
  2.010816e-013, -4.446853e-014, 2.087977e-012, 1.553871e-011,
  1.048377e-013, -3.308191e-014, 3.344774e-011, 1.713009e-010,
  2.628068e-013, -6.308238e-014, -5.74192e-011, -3.761222e-011,
  1.074936e-013, -3.543268e-014, 4.282475e-011, 1.596139e-010,
  2.070809e-013, -6.530528e-014, -3.065443e-011, 9.243863e-012,
  9.769144e-014, -4.018224e-014, 2.620641e-011, 1.345736e-010,
  1.882521e-013, -7.178902e-014, 3.342332e-012, 3.874768e-011,
  9.413038e-014, -4.762889e-014, 3.412363e-011, 1.34758e-010,
  1.814787e-013, -7.372723e-014, -3.14766e-011, -8.346501e-014,
  9.642675e-014, -5.223101e-014, 5.381179e-011, 1.263786e-010,
  1.654019e-013, -6.662643e-014, 9.716413e-012, 2.696252e-012,
  8.665091e-014, -4.538561e-014, 6.029777e-011, 1.435094e-010,
  1.636578e-013, -5.78369e-014, -2.98023e-011, 1.586713e-011,
  8.927052e-014, -3.644984e-014, 4.82045e-011, 1.526862e-010,
  1.733107e-013, -4.83922e-014, -1.656499e-013, 3.882687e-011,
  9.13648e-014, -3.134197e-014, -2.482158e-011, 9.462892e-011,
  1.664954e-013, -4.214992e-014, -4.111116e-012, 4.035602e-012,
  8.836126e-014, -2.905152e-014, 2.766406e-011, 1.104919e-010,
  1.787265e-013, -3.958536e-014, -2.912964e-011, -2.347885e-011,
  1.009842e-013, -2.824886e-014, 2.510796e-011, 1.062799e-010,
  2.014938e-013, -4.061936e-014, 6.179541e-012, -2.487077e-012,
  1.090046e-013, -2.587611e-014, 3.38128e-011, 1.354278e-010,
  1.493155e-013, -3.80877e-014, 1.113612e-011, 1.2053e-011,
  8.353005e-014, -2.453629e-014, 5.916086e-011, 1.357134e-010,
  1.449214e-013, -4.663708e-014, 2.787487e-012, 1.513175e-011,
  8.303969e-014, -3.198162e-014, 2.717526e-011, 9.442806e-011,
  1.403676e-013, -4.920768e-014, 6.691566e-012, 1.191429e-011,
  7.716222e-014, -3.447052e-014, 3.638471e-011, 1.050738e-010,
  1.169453e-013, -4.833919e-014, 2.574834e-011, 3.877486e-011,
  9.377139e-015, -2.489606e-014, 3.059893e-011, 9.254598e-011,
  1.326812e-013, -4.166396e-014, -1.976816e-012, 1.41964e-011,
  7.595768e-014, -2.99298e-014, 2.412629e-011, 9.330548e-011,
  1.305566e-013, -3.904579e-014, -1.135969e-012, 1.030366e-011,
  7.386301e-014, -2.72568e-014, 2.288575e-011, 9.191729e-011,
  1.24503e-013, -4.127687e-014, 1.66365e-012, 8.468204e-012,
  7.272412e-014, -2.792037e-014, 3.694185e-011, 9.793612e-011,
  1.226857e-013, -4.705889e-014, -2.897978e-012, 1.011207e-012,
  7.109741e-014, -3.069775e-014, 3.025728e-011, 8.274303e-011,
  1.181021e-013, -5.003852e-014, 1.886722e-011, 1.857215e-011,
  6.783025e-014, -3.454128e-014, 2.655289e-011, 7.898471e-011,
  1.128905e-013, -5.222068e-014, 1.770008e-011, 1.599726e-011,
  6.63179e-014, -3.460309e-014, 3.488202e-011, 7.784563e-011,
  8.920203e-014, -5.101494e-014, 3.643815e-012, -7.06211e-013,
  6.264197e-014, -3.767514e-014, 3.911654e-011, 7.235303e-011,
  1.149423e-013, -5.45724e-014, 7.601046e-012, 5.810469e-012,
  1.581948e-014, -2.855027e-014, 3.468298e-011, 8.105264e-011,
  1.06922e-013, -4.694195e-014, -1.195727e-012, 5.504721e-012,
  3.930034e-014, -2.971461e-014, 4.437001e-011, 7.805531e-011,
  3.688388e-014, -3.386091e-014, -8.705577e-013, 8.675368e-013,
  2.587966e-014, -2.545697e-014, 3.614879e-011, 7.21712e-011,
  8.668975e-014, -3.910718e-014, -4.202852e-012, -1.786001e-013,
  5.31488e-014, -2.949016e-014, 3.28361e-011, 7.137167e-011,
  1.225658e-013, -4.343479e-014, 5.751307e-012, 5.31898e-012,
  7.182969e-014, -2.901453e-014, 3.205417e-011, 6.402385e-011,
  1.412871e-013, -4.758028e-014, -1.696064e-011, -1.115751e-011,
  7.39097e-014, -3.088964e-014, 2.437535e-011, 5.813953e-011,
  9.172827e-014, -4.011174e-014, -6.930828e-012, -2.437087e-012,
  5.394057e-014, -2.755683e-014, 1.254107e-011, 5.159271e-011,
  8.975722e-014, -3.783008e-014, 1.867847e-011, 2.319963e-011,
  5.859022e-014, -2.53956e-014, 1.942761e-011, 5.378236e-011,
  8.637817e-014, -3.346806e-014, 1.732797e-011, 1.698543e-011,
  5.816421e-014, -2.73639e-014, 2.470183e-011, 6.611817e-011,
  8.322377e-014, -3.060738e-014, 4.0158e-011, 4.528202e-011,
  5.710474e-014, -2.391182e-014, 1.820239e-011, 6.773169e-011,
  8.527314e-014, -2.605268e-014, -8.10913e-012, 4.579385e-012,
  5.405533e-014, -1.956061e-014, -1.898929e-012, 5.151626e-011,
  8.477337e-014, -2.340227e-014, -1.671641e-011, -1.016669e-011,
  5.366791e-014, -1.450978e-014, 2.904354e-011, 6.628938e-011,
  8.074972e-014, -1.947435e-014, -1.715447e-012, -4.890975e-012,
  5.218938e-014, -1.475757e-014, 1.399673e-012, 4.645554e-011,
  1.305173e-013, -2.498884e-014, 1.012917e-011, 1.243587e-011,
  9.721048e-014, -2.105372e-014, -2.764552e-011, 2.717702e-011,
  7.911576e-014, -1.485753e-014, -2.346009e-011, -1.165992e-011,
  4.751476e-014, -1.191881e-014, 1.075811e-011, 6.53728e-011,
  7.227467e-014, -1.655657e-014, 2.528844e-011, 3.986183e-011,
  4.493182e-014, -1.050015e-014, 2.662583e-011, 7.766317e-011,
  7.447419e-014, -2.250771e-014, 1.565302e-011, 2.46517e-011,
  5.011538e-014, -1.605685e-014, 1.516512e-011, 3.802364e-011,
  6.452826e-014, -3.331452e-014, 9.031969e-013, 1.415556e-011,
  -1.100003e-014, -7.17695e-015, 2.202441e-012, 3.096485e-011,
  6.375866e-014, -3.731648e-014, 3.366114e-011, 2.163478e-011,
  2.482507e-014, -2.268155e-014, -3.098384e-011, 1.99428e-012,
  6.733179e-014, -3.662628e-014, 2.465733e-011, 4.26789e-011,
  4.550862e-014, -2.763567e-014, 1.289417e-011, 4.69977e-011,
  6.269642e-014, -3.417461e-014, 6.646818e-012, 7.838833e-012,
  4.147983e-014, -2.341609e-014, 1.185811e-011, 2.968462e-011,
  6.492892e-014, -2.72975e-014, -4.559926e-011, -3.774224e-011,
  4.19693e-014, -1.959592e-014, 6.109506e-011, 7.682138e-011,
  6.504051e-014, -2.47643e-014, -3.601787e-011, -3.302159e-011,
  4.31943e-014, -1.856481e-014, 3.361782e-011, 7.270648e-011,
  5.947212e-014, -2.539013e-014, 2.306178e-011, 4.669768e-011,
  4.094156e-014, -1.788843e-014, 1.530318e-011, 5.749476e-011,
  5.915393e-014, -2.734659e-014, 9.744009e-012, 2.673035e-011,
  3.957202e-014, -1.836521e-014, 1.161838e-011, 3.728109e-011,
  6.313176e-014, -2.760162e-014, 2.756076e-011, 2.545722e-011,
  2.715809e-014, -1.713534e-014, 4.615761e-011, 7.717046e-011,
  7.861519e-014, -3.583535e-014, 2.384383e-011, 1.357232e-011,
  -1.870095e-014, -1.359819e-014, 1.250933e-011, 3.2021e-011,
  5.292589e-014, -3.183415e-014, 6.128039e-013, -7.346434e-012,
  3.875309e-014, -2.427805e-014, 3.341035e-011, 4.897553e-011,
  5.07424e-014, -3.209079e-014, -1.384378e-011, -1.56335e-011,
  3.604935e-014, -2.567428e-014, 1.824916e-011, 3.402916e-011,
  5.063939e-014, -3.039162e-014, -1.174099e-011, -1.658486e-011,
  3.441908e-014, -2.495033e-014, 2.144797e-011, 3.804071e-011,
  1.099358e-013, -3.781102e-014, 5.181513e-012, -4.685582e-012,
  7.399414e-014, -2.862604e-014, 1.998956e-011, 3.625145e-011,
  4.938489e-014, -2.605573e-014, 8.727053e-013, -4.532307e-012,
  3.361437e-014, -2.042416e-014, 2.330671e-011, 3.99401e-011,
  4.889956e-014, -2.418711e-014, 2.963532e-011, 2.858699e-011,
  3.393512e-014, -2.005117e-014, 1.759451e-011, 1.351401e-011,
  4.561481e-014, -2.426129e-014, -2.999544e-012, 9.892144e-012,
  3.649172e-014, -2.077442e-014, 2.529079e-011, 3.792869e-011,
  4.604264e-014, -2.442882e-014, 1.517233e-011, 1.337753e-012,
  3.164577e-014, -1.861282e-014, 3.895027e-011, 5.01629e-011,
  4.596186e-014, -2.327745e-014, -8.420743e-012, 4.126429e-012,
  3.204499e-014, -1.858463e-014, 6.219204e-012, 2.915458e-011,
  4.236641e-014, -2.195009e-014, 8.629559e-012, 2.133041e-011,
  3.300284e-014, -2.098155e-014, -8.545214e-012, 6.497852e-012,
  4.431659e-014, -1.578008e-014, 6.203199e-012, -2.463553e-012,
  3.038897e-014, -1.007214e-014, -1.46834e-012, 2.41428e-011,
  4.067161e-014, -2.107379e-014, 5.060158e-011, 2.956731e-011,
  2.738708e-014, -1.057463e-014, -1.26832e-011, 1.204007e-011,
  4.311362e-014, -2.193203e-014, 5.307018e-011, 3.256881e-011,
  2.714627e-014, -1.45919e-014, 8.102672e-012, -5.122394e-014,
  4.017447e-014, -1.931558e-014, 2.51952e-011, 2.475434e-011,
  2.932443e-014, -1.621582e-014, 3.323978e-011, 3.904062e-011,
  4.023682e-014, -2.142333e-014, 8.550798e-012, 3.666661e-012,
  2.833492e-014, -2.134402e-014, 4.835024e-011, 7.112529e-011,
  4.136784e-014, -1.668328e-014, 1.217135e-011, 1.32947e-011,
  4.504403e-014, -1.502924e-014, 1.439925e-011, 2.051295e-011,
  4.949055e-014, -1.874484e-014, -2.17517e-012, -1.380997e-011,
  8.388637e-014, -2.249207e-014, 1.788443e-011, 3.237622e-011,
  3.749972e-014, -1.622372e-014, -1.539332e-011, -6.302704e-012,
  2.661774e-014, -1.569366e-014, 4.670008e-012, 1.036247e-011,
  3.474905e-014, -1.516444e-014, 3.22563e-012, 8.861174e-013,
  2.691962e-014, -1.141638e-014, 5.219898e-012, 2.788122e-011,
  3.219464e-014, -1.741825e-014, 1.230585e-011, 2.257259e-011,
  2.675842e-014, -1.156106e-014, -1.137333e-011, 1.580978e-011,
  -3.655355e-014, -7.779622e-015, 1.308307e-011, 2.5527e-012,
  2.160973e-014, -1.292996e-014, 1.102857e-011, 2.063871e-011,
  3.561718e-014, -1.455758e-014, 2.888151e-012, 4.741722e-012,
  2.388054e-014, -1.386687e-014, 2.68061e-011, 3.752298e-011,
  3.324199e-014, -1.871093e-014, 9.233744e-012, 1.403472e-011,
  2.400287e-014, -1.697681e-014, 1.767904e-011, 3.272264e-011,
  3.374721e-014, -1.820835e-014, -1.884291e-012, 5.058828e-012,
  2.366211e-014, -1.508055e-014, 3.41353e-011, 4.201361e-011,
  3.096361e-014, -1.596826e-014, 1.248335e-011, 3.783918e-012,
  2.337539e-014, -9.997171e-015, 9.656594e-013, 1.063597e-011,
  2.982508e-014, -1.708663e-014, -1.543503e-012, -1.028239e-012,
  2.151558e-014, -1.336693e-014, 1.096011e-011, 2.129836e-011,
  3.110805e-014, -1.280484e-014, 9.293609e-012, 1.019825e-011,
  2.462673e-014, -9.783448e-015, -1.057204e-011, 5.522926e-013,
  3.157295e-014, -1.557736e-014, 6.131178e-012, 2.247852e-011,
  2.202504e-014, -1.093728e-014, -3.965325e-012, 6.497816e-012,
  -1.958186e-014, -3.458062e-015, 2.248636e-011, 2.49465e-011,
  -3.328045e-015, -5.769115e-015, 1.543396e-011, 3.038676e-011,
  1.220532e-014, -8.913954e-015, 2.75086e-011, 2.435686e-011,
  1.45617e-014, -4.753092e-015, 1.174466e-011, 3.979462e-011,
  2.748624e-014, -9.516869e-015, -1.061469e-012, 1.744797e-011,
  2.230881e-014, -7.6229e-015, 4.055382e-012, 1.685172e-011,
  2.704819e-014, -9.552881e-015, -2.737878e-011, -1.817516e-011,
  2.319068e-014, -8.66499e-015, -1.044382e-012, -5.279973e-012,
  3.83982e-014, -1.668937e-014, -5.071198e-012, 1.565408e-011,
  5.038305e-014, -1.618066e-014, 4.536441e-011, 6.165136e-011,
  4.80035e-014, -1.715459e-014, 4.036882e-011, 3.945433e-011,
  5.993417e-014, -2.092737e-014, 3.72628e-011, 3.836908e-011,
  2.456417e-014, -1.418123e-014, -8.231408e-012, 6.383543e-012,
  1.701632e-014, -1.219895e-014, 5.726605e-013, 4.314221e-011,
  2.534834e-014, -1.018145e-014, 3.503814e-011, 3.423498e-011,
  1.673921e-014, -8.575894e-015, -2.036691e-013, 2.440191e-011,
  2.583052e-014, -8.833306e-015, 1.588384e-011, 1.882637e-011,
  1.725087e-014, -1.145916e-014, 7.128464e-012, 2.902741e-011,
  2.260854e-014, -1.084527e-014, 1.182349e-011, 3.097323e-012,
  2.144825e-014, -1.230251e-014, 2.403957e-011, 4.232582e-011,
  2.362078e-014, -1.379976e-014, -3.166521e-012, 1.560988e-011,
  1.918328e-014, -1.23492e-014, 1.314068e-011, 2.538285e-011,
  2.315794e-014, -1.244645e-014, -2.762254e-011, -3.939969e-012,
  2.030601e-014, -9.812682e-015, 4.288939e-012, 1.381412e-011,
  2.175615e-014, -1.559476e-014, -4.857678e-012, 1.055924e-011,
  1.680863e-014, -1.164842e-014, 3.29757e-011, 3.647747e-011,
  2.221937e-014, -1.322304e-014, -5.176497e-012, -3.691621e-012,
  8.349417e-014, -2.141058e-014, 1.252725e-011, 2.430131e-011,
  2.378043e-014, -1.431542e-014, 2.350876e-011, 2.237209e-011,
  1.647124e-014, -1.024581e-014, 3.866474e-011, 3.446857e-011,
  2.14334e-014, -1.483329e-014, 4.634492e-012, 7.287836e-012,
  1.588911e-014, -9.240925e-015, 6.047367e-012, 6.013979e-012,
  2.323357e-014, -1.339697e-014, 1.472039e-012, -1.099632e-011,
  1.783572e-014, -8.768056e-015, -2.869558e-012, 3.95481e-012,
  -3.989354e-014, -1.609991e-015, 2.313829e-011, 2.733449e-011,
  -8.439046e-016, -2.583001e-015, -2.011678e-011, 5.821551e-012,
  4.995727e-015, -7.640453e-015, 1.192894e-011, 3.215288e-011,
  1.323045e-014, -8.080452e-015, -4.940665e-012, 1.553001e-011,
  1.884724e-014, -1.065987e-014, 1.295794e-011, 5.832088e-012,
  1.43636e-014, -8.394369e-015, -9.66094e-012, 8.477203e-012,
  1.901074e-014, -1.046563e-014, -1.13692e-011, -2.141997e-012,
  1.307023e-014, -7.911823e-015, 9.103674e-012, 3.284182e-012,
  2.038497e-014, -4.312456e-015, 1.732236e-011, 1.766037e-011,
  1.458913e-014, -5.511947e-015, 7.852064e-012, 2.651743e-011,
  2.258849e-014, -5.166923e-015, -1.173092e-011, -2.19551e-011,
  1.341945e-014, -6.954103e-015, 5.002222e-012, 2.798521e-011,
  2.458813e-014, -8.005858e-015, -9.897192e-012, -1.203711e-011,
  1.62853e-014, -7.013355e-015, -7.096825e-012, -8.000235e-012,
  2.374585e-014, -3.737657e-015, -2.749826e-011, -3.28078e-011,
  1.715968e-014, -4.176409e-015, 2.808806e-011, 5.351143e-011,
  2.294741e-014, -6.856193e-015, -1.865877e-011, -1.403247e-011,
  1.799265e-014, -6.006952e-015, 3.557557e-012, 2.553756e-012,
  2.868242e-014, -5.696294e-015, 2.491844e-011, 1.959167e-011,
  2.460798e-014, -9.308517e-015, 1.904897e-011, 2.307978e-011,
  1.742935e-014, -7.959174e-015, 9.120309e-012, 3.307585e-011,
  1.208665e-014, -1.365327e-014, 1.609469e-011, 3.409033e-011,
  2.182156e-014, -1.474855e-015, 5.637348e-012, 7.15011e-012,
  1.283254e-014, -1.334033e-015, -6.740235e-011, -3.044698e-011,
  1.542714e-014, -5.528141e-015, -2.048468e-011, -7.650495e-012,
  1.770443e-014, -5.514127e-015, 2.120998e-011, 3.289527e-011,
  3.210471e-014, 1.074789e-016, 1.439945e-012, 2.497751e-012,
  2.902252e-014, 1.85603e-015, 2.954387e-013, 2.076193e-011,
  4.449299e-014, -1.212194e-015, 2.108909e-011, 1.312078e-011,
  3.136766e-014, 2.538673e-015, 2.986205e-012, 2.177358e-011,
  7.677047e-014, -4.711956e-015, -3.269529e-012, -7.066462e-012,
  4.192229e-014, -5.724014e-016, -1.629903e-012, 1.854962e-011,
  2.710956e-014, -1.801662e-015, -1.032389e-011, -1.361769e-011,
  3.046878e-014, 3.010104e-015, -1.457605e-011, -1.272825e-012,
  3.335147e-014, -1.506331e-015, -2.797718e-013, 1.636287e-012,
  3.095754e-014, -1.632992e-016, -6.566363e-012, 1.15829e-011,
  4.013393e-014, 3.109614e-015, -8.347717e-012, -6.790024e-012,
  3.144813e-014, 5.776016e-015, 4.744114e-012, 2.030539e-011,
  1.076186e-013, -6.536665e-015, 2.749495e-012, 7.163389e-012,
  5.117343e-015, 7.472398e-015, -1.226519e-012, 2.354734e-011,
  3.903701e-014, 3.359627e-015, 5.10384e-012, 7.789215e-012,
  3.285897e-014, 3.126403e-015, 6.752586e-013, 2.998738e-011,
  4.112065e-014, 2.674843e-015, 5.760883e-012, 4.032532e-012,
  3.480952e-014, 4.451057e-015, 7.964231e-013, 3.020164e-011,
  4.760619e-014, 2.230254e-014, 5.735888e-012, -1.009196e-012,
  2.892614e-014, -5.714987e-015, -7.230535e-013, 2.982319e-011,
  -1.974213e-014, 7.07803e-015, 1.303395e-011, 1.309063e-011,
  7.552196e-014, 2.242734e-015, -7.067823e-013, 2.74593e-011,
  3.662727e-014, 4.958239e-015, -2.800435e-012, -5.242297e-012,
  4.259681e-014, 3.950443e-015, -1.591235e-013, 2.968245e-011,
  3.777645e-014, 4.230011e-015, -7.786083e-012, -7.744389e-012,
  5.009011e-014, 3.286528e-015, -5.121121e-012, 2.137653e-011,
  4.43714e-014, 4.286839e-015, -2.192531e-012, 6.246917e-013,
  3.795105e-014, 2.358234e-015, -1.173613e-012, 2.333146e-011,
  4.589454e-014, 3.554519e-015, 1.547231e-012, 5.717159e-012,
  3.897096e-014, 2.96429e-015, 6.205141e-012, 3.694901e-011,
  4.961326e-014, 1.451411e-015, -2.479097e-012, -3.784171e-012,
  4.470439e-014, 4.387202e-015, 7.471007e-013, 3.240784e-011,
  4.590689e-014, 1.49457e-015, -6.62067e-012, -3.074838e-012,
  4.082735e-014, 5.795378e-015, -1.086127e-011, 1.865519e-011,
  5.05816e-014, 1.65043e-015, 1.73183e-012, 1.764823e-012,
  4.447308e-014, 4.340743e-015, -3.933152e-012, 3.128542e-011,
  5.227372e-014, 6.449083e-016, 1.725155e-013, 2.838866e-012,
  4.435403e-014, 4.439504e-015, -7.608708e-013, 3.278043e-011,
  5.428853e-014, 2.865418e-015, 1.59221e-013, 2.40762e-012,
  4.699849e-014, 8.677082e-016, -5.848229e-012, 3.229269e-011,
  5.309945e-014, -1.453465e-015, 6.975304e-013, 2.592897e-012,
  4.803798e-014, 1.018633e-016, 1.893913e-012, 3.613162e-011,
  5.434493e-014, -1.610438e-015, 2.935307e-012, 7.971616e-012,
  4.886689e-014, -1.176184e-016, 9.138359e-012, 4.443801e-011,
  5.594495e-014, -1.179588e-015, 5.697114e-012, 7.664207e-012,
  4.292999e-014, -1.775657e-016, 3.372071e-012, 3.353285e-011,
  3.746534e-014, -4.986407e-015, -3.012979e-013, -7.004891e-012,
  -1.371932e-014, 9.278864e-015, -1.957689e-012, 2.869365e-011,
  5.893358e-014, -1.366997e-014, -4.415174e-012, -6.199571e-012,
  5.788869e-014, 3.422322e-015, 1.23173e-011, 4.40114e-011,
  6.189356e-014, -1.100942e-014, -2.805194e-014, 1.43165e-012,
  5.778384e-014, 2.474983e-015, 1.196158e-013, 3.899888e-011,
  6.33735e-014, -4.990625e-015, -2.919496e-012, -6.799127e-013,
  5.796234e-014, -1.101328e-014, -5.802246e-012, 2.591834e-011,
  9.418594e-014, -1.058157e-014, 1.296516e-011, 1.398644e-011,
  1.4216e-013, -1.781168e-014, -1.15842e-011, 2.549571e-011,
  7.065912e-014, -8.326524e-015, 2.444225e-012, 1.040922e-011,
  6.59415e-014, -9.830631e-015, 1.468332e-011, 5.84985e-011,
  7.084487e-014, -8.4243e-015, -4.121117e-012, -2.003136e-012,
  6.368418e-014, -7.76837e-015, 1.13511e-011, 4.791999e-011,
  7.451902e-014, -9.162187e-015, -2.364554e-013, -1.050626e-012,
  7.07014e-014, -3.868334e-015, 7.31432e-013, 3.787099e-011,
  7.08594e-014, -8.985647e-015, 1.374492e-012, -3.182543e-011,
  7.173682e-014, -6.12774e-015, -3.640073e-012, -1.375804e-011,
  7.594504e-014, -8.150929e-015, 1.182601e-011, 1.69451e-011,
  7.267438e-014, -7.696072e-015, -3.338469e-012, 3.939207e-011,
  7.584498e-014, -5.749807e-015, 1.945276e-012, 5.126308e-012,
  8.28865e-014, -5.113182e-015, 8.539974e-012, 5.307532e-011,
  8.442579e-014, -6.917283e-015, -1.204817e-012, -5.739093e-014,
  7.685559e-014, -2.130221e-015, -7.399475e-013, 4.691915e-011,
  1.05121e-013, -1.423659e-014, 1.545486e-011, 1.276261e-011,
  8.788414e-014, -2.478111e-015, 2.738169e-013, 4.247951e-011,
  1.111672e-013, -1.61547e-014, 5.727704e-012, 6.994685e-013,
  9.122766e-014, -6.978668e-015, 7.001772e-012, 5.502513e-011,
  9.006932e-014, -1.015887e-014, 2.832452e-013, 3.236484e-012,
  8.163622e-014, -6.690687e-015, 3.194184e-012, 5.340214e-011,
  9.282574e-014, -7.929875e-015, 3.154588e-012, 4.582819e-012,
  8.772744e-014, -3.652791e-015, 2.682426e-012, 5.219007e-011,
  9.399529e-014, -4.137887e-015, 3.542152e-012, 2.09665e-012,
  7.706931e-014, 1.746888e-015, 2.344512e-012, 5.987129e-011,
  1.282914e-013, -6.337006e-015, 3.870285e-012, -5.239837e-013,
  3.334455e-014, 9.888295e-015, -2.683764e-012, 5.92852e-011,
  1.118046e-013, -6.55586e-016, -5.70917e-012, -7.677811e-012,
  9.764404e-014, 1.264635e-015, -5.379815e-012, 6.386726e-011,
  1.104617e-013, 3.665511e-016, 2.086369e-012, -5.291426e-013,
  1.014567e-013, 4.749732e-015, -3.608868e-012, 6.22494e-011,
  1.119518e-013, 1.240707e-015, -1.524007e-012, -1.056582e-012,
  1.027049e-013, 6.187472e-015, -3.361733e-012, 6.12276e-011,
  1.409534e-013, -1.256215e-015, -8.002937e-013, -1.971966e-012,
  1.828388e-013, -1.848511e-015, -6.269238e-012, 6.681754e-011,
  1.153878e-013, 6.09083e-015, -2.5951e-012, -2.914315e-012,
  1.103551e-013, 1.328239e-014, -1.486256e-011, 6.102205e-011,
  1.248294e-013, 1.198726e-014, -1.055655e-011, -1.635943e-011,
  1.172823e-013, 1.525072e-014, -5.873763e-012, 7.871011e-011,
  1.284054e-013, 1.43778e-014, 5.943318e-012, 5.269494e-012,
  1.196774e-013, 2.043664e-014, -1.27947e-011, 7.11279e-011,
  1.773076e-013, 3.265514e-014, -3.153404e-012, -1.295296e-012,
  1.144275e-013, 9.359341e-016, -6.118245e-012, 8.148051e-011,
  1.444101e-013, 2.299479e-014, -1.269585e-011, -1.83773e-011,
  1.290829e-013, 2.661193e-014, -4.741354e-012, 8.79774e-011,
  1.483353e-013, 2.736631e-014, -5.560975e-012, -5.191852e-012,
  1.351762e-013, 2.44261e-014, -1.059724e-011, 9.249945e-011,
  1.53973e-013, 1.853366e-014, 1.080347e-012, -3.57263e-013,
  1.415447e-013, 2.457276e-014, -1.464533e-011, 8.450643e-011,
  1.875701e-013, 9.437765e-015, 3.425138e-012, 1.450547e-012,
  1.182327e-013, 2.646403e-014, -1.893466e-011, 8.032831e-011,
  1.904018e-013, 1.111372e-014, 6.739418e-012, 1.144434e-011,
  1.302372e-013, 2.286519e-014, -1.691278e-011, 9.016735e-011,
  1.753331e-013, 9.705377e-015, 1.654504e-012, -1.583784e-012,
  1.590699e-013, 1.692263e-014, -1.619427e-011, 9.394272e-011,
  1.844755e-013, 5.565045e-015, 1.82191e-012, -2.807291e-012,
  1.643558e-013, 1.382323e-014, -8.635299e-012, 1.030462e-010,
  1.800278e-013, 4.983907e-015, 1.498855e-012, -5.329767e-012,
  1.896171e-013, 9.654094e-015, -1.348062e-011, 1.050452e-010,
  1.738473e-013, 4.907473e-015, 7.094448e-012, -3.519783e-013,
  2.239313e-013, 1.99215e-015, 3.046586e-012, 1.209534e-010,
  2.132952e-013, -3.731532e-015, 4.493135e-012, -4.184042e-012,
  1.839483e-013, 4.66569e-015, -1.984694e-012, 1.165734e-010,
  2.23448e-013, -9.484866e-015, 1.935969e-012, -6.204627e-012,
  1.913573e-013, 1.143041e-015, 5.734115e-013, 1.257044e-010,
  2.350736e-013, -1.504904e-014, 3.067437e-012, -4.776906e-012,
  1.983477e-013, -6.257051e-015, 6.119542e-012, 1.329204e-010,
  2.451862e-013, -1.827147e-014, 1.533282e-012, -8.22282e-012,
  2.046632e-013, -9.729357e-015, 9.356021e-012, 1.443322e-010,
  2.579276e-013, -1.888801e-014, 1.353163e-012, -7.800695e-012,
  2.154744e-013, -7.292739e-015, 6.276468e-012, 1.45402e-010,
  2.712312e-013, -1.923468e-014, 2.902622e-012, -9.999808e-012,
  2.215992e-013, -7.302645e-015, 6.140905e-012, 1.526831e-010,
  2.828809e-013, -2.198141e-014, 5.64443e-012, -9.286143e-012,
  2.282677e-013, -9.621263e-015, 6.653542e-012, 1.608474e-010,
  3.381222e-013, -3.663998e-014, 2.598205e-012, -9.993289e-012,
  2.304248e-013, -8.402614e-015, 7.671182e-013, 1.591675e-010,
  3.143628e-013, -2.628146e-014, 7.192332e-012, -1.712246e-012,
  2.442728e-013, -9.198161e-015, 3.545566e-012, 1.725731e-010,
  3.307065e-013, -2.437569e-014, 2.616834e-012, -6.898473e-012,
  2.544334e-013, -9.916546e-015, 7.308435e-012, 1.888596e-010,
  3.471444e-013, -2.092419e-014, 1.228647e-011, -1.984536e-012,
  2.617898e-013, -1.019277e-014, 4.794138e-013, 2.095197e-010,
  3.276838e-013, -1.963897e-014, 2.151527e-012, -1.552338e-011,
  2.226222e-013, 2.508644e-015, 9.903746e-012, 2.198159e-010,
  3.714321e-013, -1.9111e-014, 1.348053e-011, -5.545401e-012,
  2.658691e-013, -3.127186e-015, 3.406587e-012, 2.263552e-010,
  4.035367e-013, -2.320313e-014, 3.403941e-013, -1.644297e-011,
  2.883494e-013, -5.572078e-015, 3.001965e-013, 2.415541e-010,
  4.198863e-013, -2.745797e-014, 1.051504e-011, -9.598948e-012,
  2.955901e-013, -5.443303e-015, 3.703078e-012, 2.557368e-010,
  4.187454e-013, -2.667844e-014, 3.792013e-012, -1.496396e-011,
  3.306779e-013, -1.06613e-014, 8.701009e-012, 2.761046e-010,
  4.330193e-013, -2.409171e-014, 5.473271e-012, -9.38206e-012,
  3.521093e-013, -1.076199e-014, 8.922583e-012, 3.03073e-010,
  4.774618e-013, -1.967211e-014, 6.403096e-012, -8.421971e-012,
  3.242892e-013, 3.127299e-015, 1.220061e-012, 3.22364e-010,
  4.969565e-013, -1.197126e-014, 6.375941e-012, -8.607996e-012,
  3.378002e-013, 8.753494e-015, -3.647302e-012, 3.422512e-010,
  5.165946e-013, -1.741439e-014, 6.757891e-012, -5.280778e-012,
  3.472278e-013, 3.614448e-015, 3.021329e-012, 3.651928e-010,
  5.33785e-013, -3.023208e-014, 6.069925e-012, -2.131099e-013,
  3.569312e-013, -5.181937e-015, 5.566685e-012, 3.881915e-010,
  5.517968e-013, -4.208623e-014, 5.103875e-013, -7.493135e-013,
  3.689166e-013, -8.788979e-015, 2.526074e-011, 4.359064e-010,
  5.71024e-013, -3.657202e-014, 1.396466e-011, 2.308512e-011,
  3.847293e-013, -4.929689e-015, 2.029771e-011, 4.633018e-010,
  5.864393e-013, -2.710122e-014, -7.644679e-013, 1.135014e-011,
  4.027909e-013, 2.119577e-015, -9.350316e-012, 4.689248e-010,
  6.44995e-013, -2.712614e-014, 2.99199e-012, 1.977502e-011,
  4.153159e-013, 1.483195e-014, 9.092996e-012, 5.292107e-010,
  6.145714e-013, -2.134844e-014, 1.045259e-012, 4.401994e-011,
  4.430055e-013, 4.850742e-015, 1.290865e-011, 5.656239e-010,
  6.277688e-013, -3.434105e-014, -3.479657e-012, 5.998096e-011,
  4.679927e-013, -7.991135e-015, 1.928947e-011, 6.06873e-010,
  6.365178e-013, -3.700498e-014, 5.389416e-012, 7.617654e-011,
  5.017296e-013, -7.715074e-015, 1.050093e-011, 6.411996e-010,
  6.057265e-013, -3.605171e-014, -1.965585e-012, 9.966315e-011,
  4.857753e-013, -1.982152e-015, 1.67993e-011, 6.9528e-010,
  6.321287e-013, -4.198391e-014, 2.889151e-012, 1.287844e-010,
  5.797811e-013, -1.227558e-014, 1.280043e-011, 7.330129e-010,
  6.321898e-013, -4.770297e-014, 5.357665e-012, 1.707551e-010,
  6.463214e-013, -2.370684e-014, 3.014217e-011, 8.008906e-010,
  6.182153e-013, -5.466616e-014, 2.226174e-011, 2.239526e-010,
  7.186794e-013, -3.740589e-014, 3.175385e-011, 8.393146e-010,
  6.342083e-013, -6.772749e-014, 1.07022e-011, 2.542819e-010,
  8.422782e-013, -5.633726e-014, 4.900852e-011, 9.135284e-010,
  5.915262e-013, -5.638927e-014, 6.688409e-012, 3.134212e-010,
  9.420713e-013, -4.803577e-014, 4.618214e-011, 9.786875e-010,
  5.319893e-013, -3.945692e-014, 2.358139e-011, 3.942605e-010,
  1.060041e-012, -2.461753e-014, 2.479194e-011, 1.02986e-009,
  4.943057e-013, -2.497075e-014, 1.899333e-011, 4.586681e-010,
  1.22935e-012, -1.421811e-014, 1.948133e-011, 1.095386e-009,
  4.505828e-013, -3.076414e-014, 1.002503e-011, 5.3032e-010,
  1.442485e-012, -2.970212e-014, 4.013519e-011, 1.172181e-009,
  3.982366e-013, -4.141791e-014, 1.701139e-011, 6.287273e-010,
  1.704272e-012, -4.727431e-014, 4.220951e-011, 1.222481e-009,
  3.408969e-013, -3.854705e-014, 2.245394e-011, 7.430341e-010,
  2.024368e-012, -5.764203e-014, 4.04333e-011, 1.277768e-009,
  2.910896e-013, -2.164972e-014, 1.406265e-011, 8.611331e-010,
  2.4105e-012, -3.823311e-014, 2.684832e-011, 1.329401e-009,
  2.448071e-013, -6.199661e-015, 7.868836e-012, 9.976669e-010,
  2.881811e-012, -3.076804e-014, 2.027947e-011, 1.370699e-009,
  2.088043e-013, -3.622306e-015, 1.342833e-011, 1.146463e-009,
  3.461685e-012, -2.96563e-014, 2.010268e-011, 1.406304e-009,
  1.989464e-013, 2.855563e-014, 1.042895e-011, 1.321589e-009,
  4.16782e-012, 1.840697e-014, -5.653168e-012, 1.420966e-009,
  2.235523e-013, 6.857588e-014, -2.425847e-012, 1.503565e-009,
  5.014822e-012, 6.775032e-014, -3.314669e-011, 1.416707e-009,
  3.151031e-013, 7.443568e-014, -3.897008e-012, 1.706e-009,
  6.068935e-012, 7.091197e-014, -4.594771e-011, 1.382559e-009,
  4.563427e-013, 6.115163e-014, -7.595347e-012, 1.90863e-009,
  7.316214e-012, 3.4528e-014, -6.643561e-011, 1.306024e-009,
  7.156022e-013, 5.833215e-014, 1.054572e-011, 2.150984e-009,
  8.820429e-012, 2.054094e-014, -4.404378e-011, 1.226644e-009,
  1.229739e-012, 3.511121e-014, -2.500974e-011, 2.350879e-009,
  1.063937e-011, 6.694247e-015, -1.556845e-011, 1.084781e-009,
  1.778152e-012, 3.281757e-014, 5.351231e-013, 2.62867e-009,
  1.288441e-011, -1.444462e-014, -2.596508e-011, 8.533374e-010,
  2.698632e-012, -7.544783e-014, 3.515849e-011, 2.880592e-009,
  1.556118e-011, -1.450015e-013, 1.872696e-011, 5.798804e-010,
  4.007611e-012, -2.442058e-013, 7.499283e-011, 3.098898e-009,
  1.878897e-011, -3.388591e-013, 8.027488e-011, 2.083976e-010,
  5.837667e-012, -2.812011e-013, 7.867215e-011, 3.29154e-009,
  2.2648e-011, -3.609682e-013, 4.133007e-011, -3.402156e-010,
  8.395165e-012, -3.394394e-013, 8.070093e-011, 3.430367e-009,
  2.731593e-011, -3.79416e-013, 3.590155e-011, -9.770327e-010,
  1.191272e-011, -5.548338e-013, 9.947956e-011, 3.465505e-009,
  3.287838e-011, -5.356333e-013, 6.121403e-011, -1.788764e-009,
  1.675033e-011, -9.940949e-013, 1.512652e-010, 3.346268e-009,
  3.963828e-011, -8.487225e-013, 1.113552e-010, -2.837146e-009,
  2.331374e-011, -1.494329e-012, 1.993057e-010, 3.018295e-009,
  4.77331e-011, -1.14569e-012, 1.489672e-010, -4.156047e-009,
  3.22682e-011, -2.194283e-012, 2.619639e-010, 2.364115e-009,
  5.761127e-011, -1.474765e-012, 1.811586e-010, -5.830743e-009,
  4.447068e-011, -2.888022e-012, 2.868931e-010, 1.220303e-009,
  6.960608e-011, -1.665043e-012, 2.178588e-010, -7.910629e-009,
  6.132416e-011, -4.510241e-012, 4.160805e-010, -5.523529e-010,
  8.414874e-011, -2.256195e-012, 3.055668e-010, -1.050987e-008,
  8.434614e-011, -6.652011e-012, 5.474788e-010, -3.260096e-009,
  1.017015e-010, -2.925227e-012, 4.001992e-010, -1.370136e-008,
  1.160503e-010, -8.032507e-012, 5.251358e-010, -7.317548e-009,
  1.214451e-010, -3.234236e-012, 3.631795e-010, -1.772033e-008,
  1.618338e-010, -1.024138e-011, 5.611408e-010, -1.342293e-008,
  1.497695e-010, -3.348501e-012, 4.191002e-010, -2.270524e-008,
  2.277146e-010, -1.503343e-011, 7.482155e-010, -2.266895e-008,
  1.814005e-010, -3.606599e-012, 5.934684e-010, -2.909649e-008,
  3.243358e-010, -1.936742e-011, 8.687021e-010, -3.681619e-008,
  2.234989e-010, -3.631013e-012, 7.142614e-010, -3.724034e-008,
  4.699615e-010, -2.413357e-011, 9.13483e-010, -5.848291e-008,
  2.764702e-010, -3.280209e-012, 7.850568e-010, -4.758879e-008,
  7.033836e-010, -2.982035e-011, 1.088961e-009, -9.34023e-008,
  3.464365e-010, -2.379531e-012, 9.317757e-010, -6.126938e-008,
  1.0934e-009, -3.614949e-011, 1.895498e-009, -1.51362e-007,
  4.403224e-010, -5.308558e-015, 1.385896e-009, -7.948571e-008,
  1.788187e-009, -5.71705e-011, 5.059508e-009, -2.568679e-007,
  5.677013e-010, 4.388964e-012, 2.646505e-009, -1.05033e-007,
  3.021074e-009, -1.114167e-010, 1.340282e-008, -4.700845e-007,
  7.4031e-010, 9.883075e-012, 5.008622e-009, -1.42433e-007,
  4.193214e-009, -2.673306e-010, 3.801919e-008, -9.731331e-007,
  9.018332e-010, 1.804496e-011, 9.285746e-009, -2.011918e-007,
  -9.427018e-010, -5.703445e-010, 1.065592e-007, -2.154999e-006,
  8.354279e-010, 2.801384e-011, 1.671026e-008, -2.842552e-007,
  -1.071026e-008, -6.001083e-010, 1.676836e-007, -3.546997e-006,
  8.758912e-010, 3.746842e-011, 1.991678e-008, -3.466794e-007,
  -1.271318e-008, -5.952103e-010, 1.66654e-007, -3.960506e-006,
  9.349967e-010, 2.213906e-011, 1.676077e-008, -3.579669e-007,
  -9.71813e-009, -1.015579e-009, 1.13272e-007, -3.337185e-006,
  1.033134e-009, -1.100814e-011, 1.160062e-008, -3.111199e-007,
  4.886281e-010, -1.093377e-009, 4.804146e-008, -1.914745e-006,
  1.102517e-009, -7.239995e-012, 7.655689e-009, -2.305511e-007,
  4.25131e-009, -4.390649e-010, 1.769257e-008, -8.657223e-007,
  8.76643e-010, 4.639314e-012, 4.819003e-009, -1.708782e-007,
  2.869743e-009, -9.20149e-011, 6.156081e-009, -4.28977e-007,
  6.82321e-010, 5.267318e-012, 2.347915e-009, -1.278656e-007,
  1.693569e-009, -1.624921e-011, 1.721391e-009, -2.399067e-007,
  5.304592e-010, 1.281146e-012, 9.452167e-010, -9.74172e-008,
  1.040998e-009, -2.037622e-011, 8.352111e-010, -1.437079e-007,
  4.15202e-010, -2.21928e-012, 6.355179e-010, -7.503391e-008,
  6.765284e-010, -2.667117e-011, 8.343353e-010, -9.00898e-008,
  3.306696e-010, -4.960928e-012, 6.720416e-010, -5.868834e-008,
  4.581403e-010, -3.081656e-011, 1.260704e-009, -5.78505e-008,
  2.668947e-010, -6.396909e-012, 9.649074e-010, -4.633769e-008,
  3.18531e-010, -2.471369e-011, 1.335894e-009, -3.738214e-008,
  2.173339e-010, -5.766553e-012, 9.900825e-010, -3.673541e-008,
  2.263841e-010, -1.584318e-011, 1.13221e-009, -2.396904e-008,
  1.787702e-010, -4.243623e-012, 8.419744e-010, -2.923567e-008,
  1.634353e-010, -8.648461e-012, 8.335717e-010, -1.489205e-008,
  1.475234e-010, -2.755724e-012, 6.102803e-010, -2.326084e-008,
  1.189527e-010, -7.284178e-012, 8.141285e-010, -8.779125e-009,
  1.22366e-010, -2.89029e-012, 6.269187e-010, -1.844328e-008,
  8.711883e-011, -5.669668e-012, 7.795317e-010, -4.671155e-009,
  1.027987e-010, -2.399929e-012, 6.574964e-010, -1.456411e-008,
  6.406466e-011, -4.964766e-012, 7.390972e-010, -1.876957e-009,
  8.569561e-011, -2.325884e-012, 6.654038e-010, -1.142886e-008,
  4.719649e-011, -3.592363e-012, 5.968701e-010, 1.754851e-011,
  7.150928e-011, -1.752856e-012, 5.740942e-010, -8.870981e-009,
  3.465017e-011, -1.789226e-012, 3.708126e-010, 1.293953e-009,
  5.969047e-011, -7.569419e-013, 4.020063e-010, -6.78656e-009,
  2.540844e-011, -1.286347e-013, 1.447579e-010, 2.124606e-009,
  4.980082e-011, 1.843007e-013, 2.203365e-010, -5.054758e-009,
  1.851498e-011, -1.087594e-013, 1.269489e-010, 2.611084e-009,
  4.154966e-011, 6.242663e-014, 1.883372e-010, -3.683723e-009,
  1.337921e-011, -4.309588e-013, 1.570511e-010, 2.877105e-009,
  3.468285e-011, -2.04184e-013, 2.180725e-010, -2.557705e-009,
  9.563634e-012, -2.909068e-013, 8.704242e-011, 2.942862e-009,
  2.899522e-011, -9.135027e-014, 1.495038e-010, -1.671632e-009,
  6.795568e-012, -1.024072e-013, 5.52366e-011, 2.924325e-009,
  2.428965e-011, 7.414758e-014, 1.195815e-010, -9.362269e-010,
  4.742986e-012, -2.529338e-014, -1.984073e-012, 2.784008e-009,
  2.03165e-011, 1.112957e-013, 7.107855e-011, -3.903489e-010,
  3.248418e-012, -7.738958e-014, 3.062265e-011, 2.670832e-009,
  1.708553e-011, 2.431099e-014, 8.976604e-011, 3.863133e-011,
  2.202645e-012, -6.225549e-014, 3.555036e-011, 2.51363e-009,
  1.42621e-011, 1.309743e-014, 6.769914e-011, 3.787409e-010,
  1.451111e-012, -2.103056e-014, -9.699279e-013, 2.305435e-009,
  1.198526e-011, 5.863775e-014, 3.592195e-011, 6.416704e-010,
  9.150556e-013, 3.043378e-014, -5.4129e-012, 2.115577e-009,
  1.003701e-011, 1.035088e-013, 1.832022e-011, 8.439494e-010,
  5.618207e-013, 1.55837e-014, -1.896909e-012, 1.934085e-009,
  8.430762e-012, 7.11348e-014, 1.666689e-011, 9.969077e-010,
  3.288901e-013, -4.263097e-015, 1.330934e-011, 1.751007e-009,
  7.092786e-012, 2.78422e-014, 2.720496e-011, 1.10293e-009,
  1.942239e-013, -2.343375e-014, 1.416681e-011, 1.560714e-009,
  5.956754e-012, 1.043197e-015, 3.254549e-011, 1.151714e-009,
  1.233169e-013, -3.407748e-014, 3.023215e-011, 1.41171e-009,
  5.009377e-012, -3.233923e-014, 2.873671e-011, 1.185925e-009,
  9.546746e-014, -1.94857e-014, -2.541743e-012, 1.225736e-009,
  4.219055e-012, 1.010258e-014, 3.914567e-012, 1.197546e-009,
  9.922696e-014, 3.130716e-014, -1.951524e-011, 1.084118e-009,
  3.554308e-012, 9.62522e-014, -4.664377e-011, 1.187791e-009,
  1.223784e-013, 4.862298e-014, -9.624818e-012, 9.576457e-010,
  2.999179e-012, 1.325139e-013, -6.132805e-011, 1.177265e-009,
  1.647204e-013, 5.010548e-014, -1.500654e-011, 8.395983e-010,
  2.532585e-012, 1.135152e-013, -4.591893e-011, 1.164561e-009,
  2.104442e-013, 2.352477e-014, -1.260555e-011, 7.310582e-010,
  2.146994e-012, 5.563706e-014, -1.735229e-011, 1.131294e-009,
  2.605059e-013, -2.836906e-014, 4.011713e-012, 6.518934e-010,
  1.82739e-012, -5.031097e-014, 3.812558e-011, 1.08953e-009,
  3.075035e-013, -7.065082e-014, 2.952562e-011, 5.774194e-010,
  1.557228e-012, -1.114167e-013, 7.8358e-011, 1.03433e-009,
  3.478198e-013, -5.938339e-014, 3.345224e-011, 4.929059e-010,
  1.342737e-012, -9.713433e-014, 8.93062e-011, 1.012254e-009,
  3.928056e-013, -3.436623e-014, 1.607371e-011, 4.10709e-010,
  1.159179e-012, -6.11515e-014, 3.409993e-011, 9.326075e-010,
  4.525712e-013, -2.089615e-014, 1.289558e-011, 3.610688e-010,
  9.751377e-013, -1.475592e-014, 1.841442e-011, 8.941082e-010,
  4.574403e-013, 2.217468e-015, -1.735194e-011, 2.829411e-010,
  8.860299e-013, 5.355624e-015, 2.576981e-011, 8.778328e-010,
  4.859053e-013, 1.386964e-014, -8.270087e-012, 2.480308e-010,
  7.820175e-013, 7.52103e-015, -5.612917e-013, 8.183796e-010,
  5.050334e-013, 6.1135e-016, -6.864827e-013, 2.156932e-010,
  6.948992e-013, -3.189187e-015, 2.623208e-011, 7.835317e-010,
  4.647788e-013, 1.097299e-016, 3.347566e-012, 1.770203e-010,
  6.105166e-013, -2.659193e-014, 2.406534e-011, 7.219714e-010,
  5.265479e-013, -3.560652e-014, -1.127601e-011, 1.259641e-010,
  5.687384e-013, -4.805435e-014, 3.546159e-011, 6.669062e-010,
  5.423556e-013, -4.6116e-014, -9.214469e-012, 1.084626e-010,
  5.245468e-013, -6.349615e-014, 5.584556e-011, 6.443144e-010,
  5.417057e-013, -5.569583e-014, 3.781351e-012, 1.051511e-010,
  4.84831e-013, -7.187058e-014, 7.196373e-011, 6.218642e-010,
  5.873224e-013, -7.549726e-014, -3.842855e-012, 7.504858e-011,
  4.622642e-013, -8.55171e-014, 5.640943e-011, 5.564832e-010,
  5.628092e-013, -7.685656e-014, 4.8602e-012, 6.046061e-011,
  4.169763e-013, -7.917957e-014, 5.943538e-011, 5.303898e-010,
  5.262653e-013, -7.386102e-014, -4.663549e-012, 3.927699e-011,
  3.994318e-013, -7.702224e-014, 7.731783e-011, 5.133352e-010,
  5.2436e-013, -7.150304e-014, -2.980299e-011, 3.083228e-012,
  3.775715e-013, -6.577315e-014, 5.901262e-011, 4.680111e-010,
  5.137432e-013, -5.329159e-014, -5.716701e-012, 8.767201e-012,
  3.677717e-013, -5.583989e-014, 4.163149e-011, 4.348281e-010,
  5.022107e-013, -3.539317e-014, -1.363719e-011, -1.333997e-011,
  3.473851e-013, -2.812211e-014, 4.007509e-011, 4.278143e-010,
  4.928966e-013, -1.560745e-014, -1.090584e-011, 2.094003e-012,
  3.382685e-013, -2.381105e-014, 1.320706e-011, 3.771454e-010,
  4.836462e-013, -1.606096e-014, -1.502218e-011, -1.155733e-011,
  3.296538e-013, -2.121987e-014, 2.206968e-011, 3.762818e-010,
  4.663376e-013, -2.556374e-014, -1.583429e-011, -1.990621e-011,
  3.078974e-013, -2.545162e-014, 3.471719e-011, 3.752999e-010,
  4.85328e-013, -6.050178e-014, -1.557271e-011, -2.025814e-011,
  2.66779e-013, -4.865974e-014, 4.543832e-011, 3.296002e-010,
  4.389392e-013, -7.480934e-014, 1.545856e-011, -4.017528e-012,
  2.896047e-013, -6.659451e-014, 4.837274e-011, 2.874397e-010,
  4.175354e-013, -8.796121e-014, -2.364131e-011, -3.244504e-011,
  2.834255e-013, -7.606711e-014, 5.915455e-011, 2.721193e-010,
  4.001553e-013, -9.873245e-014, 1.661402e-011, 4.351955e-012,
  2.746469e-013, -8.563062e-014, 6.730645e-011, 2.678811e-010,
  3.21913e-013, -9.417497e-014, -1.296345e-012, -9.594861e-012,
  2.46975e-013, -9.118891e-014, 5.541901e-011, 2.355173e-010,
  3.67717e-013, -1.137076e-013, 1.150019e-011, 5.95758e-012,
  2.567837e-013, -1.048524e-013, 6.692467e-011, 2.278589e-010,
  3.518609e-013, -1.111587e-013, 9.973486e-012, -6.823062e-012,
  2.519404e-013, -1.009806e-013, 4.777545e-011, 1.911853e-010,
  3.4183e-013, -8.581064e-014, 9.499877e-012, -2.713518e-012,
  2.417488e-013, -7.384836e-014, 6.138111e-011, 2.262843e-010,
  3.85116e-013, -6.800172e-014, 1.42979e-011, 1.483954e-012,
  2.395155e-013, -5.585381e-014, 4.136347e-011, 2.046711e-010,
  3.330889e-013, -5.508421e-014, 2.811261e-012, -1.601262e-011,
  2.319217e-013, -4.04985e-014, 3.069013e-011, 1.817685e-010,
  3.007427e-013, -5.328621e-014, -4.644762e-012, -2.242481e-011,
  2.26101e-013, -4.227388e-014, 3.196075e-011, 1.803019e-010,
  2.876252e-013, -5.357585e-014, 1.458697e-012, -1.869202e-011,
  2.176211e-013, -4.138396e-014, 3.015626e-011, 1.651489e-010,
  2.747872e-013, -4.700002e-014, 4.666776e-012, -9.395911e-012,
  2.091624e-013, -3.924594e-014, 1.869661e-011, 1.423366e-010,
  2.64671e-013, -4.080281e-014, 3.505818e-012, -5.185456e-012,
  2.010934e-013, -4.03339e-014, 1.785086e-011, 1.350741e-010,
  2.533036e-013, -3.850619e-014, -2.267214e-012, -1.771956e-011,
  1.958857e-013, -4.188267e-014, 2.680948e-011, 1.435593e-010,
  2.408758e-013, -4.62595e-014, -8.072997e-012, -1.953772e-011,
  1.887077e-013, -4.453289e-014, 9.638151e-012, 1.158934e-010,
  2.385133e-013, -3.861403e-014, 2.011401e-011, 8.900666e-012,
  1.770613e-013, -3.364112e-014, 1.448814e-011, 1.218926e-010,
  2.48403e-013, -3.615041e-014, 1.42081e-011, 9.850502e-012,
  1.457668e-013, -2.848448e-014, 7.907993e-012, 1.112627e-010,
  2.118278e-013, -2.040422e-014, -1.161218e-011, -1.66426e-011,
  1.731698e-013, -3.11201e-014, 1.909448e-011, 1.114178e-010,
  2.045158e-013, -2.567039e-014, 1.534123e-011, 1.540404e-011,
  1.702282e-013, -1.900542e-014, 3.318661e-011, 1.365142e-010,
  1.966342e-013, -2.630213e-014, -4.78322e-012, 2.218091e-012,
  1.644016e-013, -1.77152e-014, 8.054763e-012, 1.029674e-010,
  1.225243e-013, -1.498037e-014, -5.829578e-012, -2.764948e-012,
  1.363728e-013, -1.305162e-014, -5.097374e-011, 4.751409e-011,
  1.806869e-013, -2.322323e-014, 1.621535e-011, 1.35882e-011,
  1.505666e-013, -2.252671e-014, 1.810854e-011, 9.512995e-011,
  1.763312e-013, -4.010702e-014, 5.886684e-012, 4.429131e-012,
  1.519874e-013, -3.100998e-014, 6.65169e-012, 7.112113e-011,
  1.679788e-013, -3.708706e-014, 3.434854e-012, 2.293502e-011,
  1.392448e-013, -4.305018e-014, -1.831257e-011, 6.837732e-011,
  2.271723e-013, -5.134593e-014, 2.398575e-011, 3.44974e-012,
  1.43251e-013, -4.306351e-014, -1.124743e-011, 7.334864e-011,
  1.659783e-013, -4.380496e-014, -8.312348e-012, -2.012498e-011,
  1.350935e-013, -4.241298e-014, 4.541993e-012, 4.894534e-011,
  1.47508e-013, -4.45493e-014, -1.669241e-011, -2.542729e-011,
  1.327648e-013, -5.551689e-014, 2.569311e-011, 8.506597e-011,
  1.37086e-013, -5.805575e-014, -2.036245e-011, -4.423557e-011,
  1.298439e-013, -4.443715e-014, 2.010201e-011, 5.909193e-011,
  1.358368e-013, -5.53294e-014, -3.852649e-011, -5.304615e-011,
  9.284239e-014, -4.243086e-014, 2.403085e-011, 7.320779e-011,
  1.336476e-013, -4.164333e-014, -9.097682e-013, 6.400184e-014,
  1.024452e-013, -3.754524e-014, 1.882581e-011, 5.718203e-011,
  1.282341e-013, -1.635031e-014, -3.976113e-011, -1.289343e-011,
  1.166621e-013, -3.693441e-014, 1.347076e-011, 7.922524e-011,
  1.272416e-013, -2.270625e-014, -1.49689e-012, 9.883178e-012,
  1.122435e-013, -2.240784e-014, -1.491528e-011, 3.152971e-011,
  9.957562e-014, -2.583595e-014, -4.093942e-012, -7.839784e-012,
  1.138396e-013, -3.215423e-014, 1.545562e-011, 5.160043e-011,
  6.361991e-014, -1.40328e-014, -2.636598e-012, -5.08373e-012,
  1.176672e-013, -2.486271e-014, 3.555073e-011, 8.337092e-011,
  1.102413e-013, -2.446321e-014, -3.070406e-012, -1.359492e-011,
  1.085274e-013, -2.527632e-014, 4.139499e-012, 4.660251e-011,
  1.031379e-013, -2.812049e-014, -1.17526e-011, 1.795614e-012,
  9.619433e-014, -2.891532e-014, 1.662547e-011, 5.343917e-011,
  1.014884e-013, -3.711752e-014, -7.620782e-012, -3.993177e-012,
  9.257852e-014, -3.520442e-014, 2.390201e-011, 7.140319e-011,
  1.299747e-013, -4.003689e-014, -1.920473e-011, -1.952955e-011,
  1.506522e-013, -4.269169e-014, 3.438147e-011, 7.747376e-011,
  9.008275e-014, -3.270018e-014, 1.446495e-012, 4.925016e-012,
  8.726105e-014, -3.369224e-014, 1.443794e-011, 5.864374e-011,
  9.015787e-014, -2.873586e-014, 1.571684e-011, 1.360137e-011,
  8.472026e-014, -2.346815e-014, 1.468729e-011, 4.905411e-011,
  8.791191e-014, -2.732054e-014, 1.404563e-011, 4.191072e-012,
  8.075606e-014, -2.66792e-014, 1.828209e-011, 6.035367e-011,
  8.681256e-014, -3.200876e-014, 2.855349e-011, 3.316343e-011,
  7.905627e-014, -2.517158e-014, 9.002669e-012, 3.569252e-011,
  8.128693e-014, -3.221815e-014, 6.049167e-012, 9.968464e-012,
  7.649378e-014, -2.869662e-014, 2.090464e-011, 4.23224e-011,
  7.912791e-014, -3.871003e-014, 1.018719e-011, 4.50728e-012,
  7.542219e-014, -3.446761e-014, 4.056103e-011, 6.392794e-011,
  1.035388e-013, -4.378238e-014, -7.502029e-012, -1.110501e-011,
  6.101119e-014, -3.257413e-014, 4.116816e-011, 6.285025e-011,
  4.041567e-014, -2.512159e-014, -7.926584e-013, -1.486842e-011,
  3.680051e-014, -2.768699e-014, 2.435247e-011, 4.785406e-011,
  5.14776e-014, -3.065902e-014, 1.21589e-011, 1.527201e-011,
  5.304299e-014, -3.136457e-014, 5.117741e-012, 1.828313e-011,
  1.130161e-014, -1.235056e-014, 2.437153e-011, 3.850115e-011,
  7.219172e-014, -2.931046e-014, 3.310449e-011, 5.737318e-011,
  5.64544e-014, -3.073954e-014, 1.944916e-011, 2.309595e-011,
  6.970032e-014, -2.894112e-014, 1.685796e-011, 3.877576e-011,
  8.87132e-014, -3.146977e-014, 6.580968e-012, 1.861167e-011,
  7.856975e-014, -3.120973e-014, 3.062724e-011, 5.433519e-011,
  1.111772e-013, -3.708421e-014, 3.737119e-012, 6.403904e-013,
  8.741536e-014, -2.901232e-014, 1.376055e-011, 3.272357e-011,
  5.993154e-014, -2.655642e-014, 2.973303e-011, 1.935446e-011,
  6.177962e-014, -2.101497e-014, 9.172304e-012, 3.308698e-011,
  6.188275e-014, -2.995342e-014, -1.886567e-012, -5.876419e-012,
  6.066128e-014, -2.44189e-014, 2.230877e-011, 4.16264e-011,
  6.01868e-014, -2.621429e-014, 4.294975e-012, 1.466707e-011,
  5.65332e-014, -2.560368e-014, 2.879224e-011, 4.200709e-011,
  5.659995e-014, -2.60946e-014, -4.531499e-013, 6.718661e-012,
  5.347988e-014, -2.277638e-014, 1.646542e-011, 4.379913e-011,
  6.39877e-014, -1.737872e-014, -2.662387e-012, 5.883182e-012,
  5.219184e-014, -2.135397e-014, -1.492705e-011, 2.060904e-011,
  5.790895e-014, -1.05187e-014, -1.973602e-011, -1.374881e-011,
  5.420564e-014, -1.474234e-014, 1.162351e-011, 3.525318e-011,
  5.409155e-014, -1.121899e-014, -1.647639e-011, -7.574663e-012,
  5.887991e-014, -1.495925e-014, 1.979901e-011, 4.106393e-011,
  -1.479883e-014, -2.350135e-015, 2.491114e-012, 1.144885e-011,
  3.579845e-014, -1.346102e-014, 1.72172e-011, 3.44263e-011,
  5.183189e-014, -1.064563e-014, -4.073459e-011, -4.276663e-011,
  5.186466e-014, -1.169954e-014, -1.386874e-011, 2.039414e-011,
  4.497379e-014, -1.065401e-014, 3.535859e-012, 1.361558e-011,
  4.52855e-014, -2.229114e-014, 2.372795e-012, 1.113256e-011,
  4.727865e-014, -2.564601e-014, -1.116999e-011, -5.507716e-013,
  4.929296e-014, -1.755267e-014, -5.09078e-012, -1.01891e-011,
  6.106855e-014, -2.314081e-014, 9.568303e-012, -1.088666e-011,
  1.09173e-013, -1.941779e-014, 9.386161e-012, 5.248973e-011,
  5.704932e-014, -2.383768e-014, -4.452127e-011, -4.399959e-011,
  5.966342e-014, -1.784139e-014, 1.829872e-011, 4.847606e-011,
  3.543166e-014, -2.235065e-014, -3.279192e-012, -1.070538e-011,
  4.739446e-014, -1.576845e-014, 3.620532e-011, 4.246379e-011,
  4.45312e-014, -2.574455e-014, -2.562524e-011, -2.175455e-011,
  4.709374e-014, -1.831894e-014, 2.46496e-011, 3.042613e-011,
  3.691838e-014, -1.682255e-014, -1.698751e-011, -2.619685e-011,
  4.794356e-014, -1.624893e-014, 3.69927e-011, 4.770669e-011,
  4.236355e-014, -1.185511e-014, 4.280844e-011, 2.040556e-011,
  4.277353e-014, -1.426776e-014, 1.352059e-011, 2.777285e-011,
  3.873145e-014, -2.556247e-014, 1.651299e-011, 3.079529e-012,
  3.936679e-014, -2.059702e-014, 2.985179e-011, 2.239401e-011,
  4.032729e-014, -1.785321e-014, 1.295589e-012, -2.466157e-012,
  3.641321e-014, -1.917134e-014, 1.007682e-011, 2.464418e-011,
  3.572087e-014, -1.823904e-014, -1.904205e-011, -9.172493e-012,
  2.185765e-014, -2.355885e-014, 1.260331e-011, 2.316314e-011,
  1.466543e-014, -2.018372e-014, -1.328948e-011, -2.979388e-012,
  -2.435614e-014, -2.007185e-014, 2.392692e-011, 2.778906e-011,
  3.737295e-014, -2.541227e-014, 1.049262e-012, 4.924149e-013,
  3.262591e-014, -2.071119e-014, 8.373055e-012, 8.975498e-012,
  3.637656e-014, -2.443751e-014, 1.098553e-011, 5.877747e-012,
  3.275107e-014, -1.637736e-014, 1.274886e-011, 1.300406e-011,
  3.711643e-014, -1.870837e-014, -1.758713e-012, -4.545495e-012,
  3.651141e-014, -1.707223e-014, 1.553356e-011, 3.580475e-011,
  7.356943e-014, -3.161061e-014, -1.854186e-011, -2.422656e-011,
  8.95008e-014, -2.191071e-014, 1.711446e-011, 1.616918e-011,
  3.370832e-014, -2.150688e-014, -2.520532e-011, -2.014948e-011,
  3.299325e-014, -1.920854e-014, 1.159195e-011, 8.584029e-012,
  3.399065e-014, -8.384222e-015, -2.093212e-011, -1.83396e-011,
  3.59355e-014, -1.143566e-014, 7.531755e-012, 2.295149e-011,
  3.206145e-014, -9.082762e-015, -1.449016e-011, -2.029787e-011,
  3.575659e-014, -7.801134e-015, 1.661968e-011, 7.618707e-012,
  2.641693e-014, -7.59151e-015, -9.253682e-012, -1.750549e-011,
  3.012114e-014, -1.805491e-014, 3.330001e-011, 4.52694e-011,
  3.503805e-014, -2.255616e-014, 2.352501e-011, 3.101908e-011,
  2.04573e-014, -1.825755e-014, 1.953061e-011, 1.425391e-011,
  3.118458e-014, -2.90556e-014, -1.341251e-011, -9.053781e-012,
  3.032232e-014, -1.591157e-014, 2.559117e-011, 2.655985e-011,
  3.245039e-014, -1.221482e-014, -8.947623e-012, -2.87807e-011,
  3.227614e-014, -5.864203e-015, 3.180622e-012, 2.626794e-011,
  3.231126e-014, -8.517761e-015, -2.48567e-012, -7.87683e-012,
  3.2914e-014, -1.092993e-014, -6.586654e-012, 1.56505e-011,
  2.877605e-014, -1.866265e-014, -1.079315e-011, -1.479386e-011,
  2.843647e-014, -1.490937e-014, -3.327958e-011, -9.231115e-012,
  2.991085e-014, -2.180908e-014, -5.511674e-012, -5.198121e-012,
  3.458497e-014, -1.261733e-014, -3.268871e-011, -2.263487e-011,
  2.337698e-014, -1.893308e-014, -1.173905e-011, -1.760915e-011,
  2.31839e-014, -2.164961e-014, -1.147382e-012, 4.310043e-012,
  1.742573e-014, -1.175334e-014, 4.51716e-012, 2.940899e-014,
  6.237377e-015, -1.194284e-014, 3.07928e-011, 1.906511e-011,
  1.944051e-015, -2.533462e-015, 1.89667e-011, 6.924823e-012,
  -2.545529e-014, -6.679589e-016, 2.451186e-011, 2.946178e-011,
  3.030308e-014, -9.73481e-015, -1.012134e-011, -2.016626e-012,
  2.897791e-014, -9.047961e-015, 2.962317e-011, 6.409014e-011,
  2.536384e-014, -1.772438e-014, -8.206978e-012, -2.233003e-011,
  2.955534e-014, -1.575971e-014, 6.751075e-012, 1.846967e-011,
  2.787277e-014, -1.274871e-014, -3.888999e-011, -2.111129e-011,
  2.372545e-014, -1.233767e-014, -8.149763e-012, 1.42054e-012,
  6.457947e-014, -2.567262e-014, 5.048067e-012, 7.270087e-012,
  7.903549e-014, -2.248442e-014, -2.917023e-012, 8.261616e-012,
  2.370654e-014, -1.439824e-014, -1.365167e-011, -5.80732e-012,
  1.970018e-014, -1.298058e-014, 2.397923e-012, 1.404686e-011,
  2.332345e-014, -1.703231e-014, 1.197289e-011, 9.626902e-012,
  2.016106e-014, -1.387635e-014, 3.03548e-011, 3.920929e-011,
  2.442523e-014, -7.61968e-015, -8.254354e-012, -1.570343e-011,
  2.272003e-014, -9.266235e-015, 1.06628e-011, 2.621106e-011,
  2.040801e-014, -9.395378e-015, -2.226852e-011, -1.124933e-011,
  2.040999e-014, -8.978802e-015, -3.868151e-012, -3.347254e-012,
  2.013337e-014, -1.086828e-014, 2.121921e-011, 2.83113e-011,
  2.126717e-014, -1.164537e-014, 4.943668e-012, -3.29734e-012,
  1.635308e-014, -1.071882e-014, 8.200361e-012, -2.075307e-012,
  2.19546e-014, -9.368487e-015, 2.012947e-011, 3.480838e-011,
  2.230688e-014, -1.073173e-014, -1.868463e-011, -3.415356e-012,
  2.111297e-014, -5.298187e-015, -2.149826e-011, -6.640598e-012,
  -1.393283e-014, -7.369963e-015, -1.769509e-011, -3.151789e-011,
  -1.719066e-014, -3.243075e-015, 9.254543e-012, 2.001534e-011,
  5.727744e-015, -1.28728e-014, -7.65938e-013, -2.502423e-012,
  5.171967e-015, -4.229476e-015, 1.474116e-011, 2.208438e-011,
  1.712095e-014, -1.176248e-014, -3.405699e-011, -2.908328e-011,
  1.435823e-014, -9.629767e-015, 3.020234e-011, 2.637003e-011,
  1.727751e-014, -1.137117e-015, -2.110535e-011, -1.761491e-011,
  1.620711e-014, -1.581447e-015, -4.832732e-013, -3.921226e-012,
  7.425214e-015, -1.328608e-014, -1.058723e-011, 3.273327e-012,
  4.438524e-014, -6.561734e-015, 8.921603e-012, 1.487786e-011,
  1.847743e-015, -8.209237e-015, -2.94708e-011, -9.335731e-012,
  6.756595e-014, -1.859735e-014, 1.641462e-012, 8.53262e-012,
  1.676694e-014, 1.015009e-015, 1.332749e-011, 2.505081e-011,
  2.112122e-014, -1.092598e-014, 3.359229e-011, 3.612526e-011,
  1.990238e-014, 3.06466e-016, 1.355694e-011, 1.858854e-011,
  2.687211e-014, -8.742673e-016, 3.170282e-012, 1.522659e-011,
  1.329547e-014, -1.865974e-014, 1.995079e-011, 6.694581e-012,
  2.135847e-014, -6.26157e-015, 3.043433e-011, 1.210889e-011,
  1.109414e-014, -7.392251e-015, 1.879959e-012, 1.470208e-011,
  1.680948e-014, -8.759332e-015, -7.9912e-012, 4.256343e-012,
  1.673796e-014, -5.7915e-015, -9.968631e-012, -1.011046e-011,
  1.916721e-014, -7.094924e-015, -2.487469e-013, 2.049145e-011,
  1.454878e-014, -1.464186e-014, -3.47083e-012, 7.215093e-012,
  1.790831e-014, -8.466575e-015, 6.733714e-012, 1.595988e-011,
  2.654085e-014, -7.576057e-015, -1.96598e-011, -7.669107e-012,
  1.84834e-014, -8.151381e-015, 1.261334e-011, -1.805365e-012,
  3.080037e-014, -1.535259e-014, 2.341047e-012, 2.534148e-011,
  -4.961856e-014, 6.815992e-015, -7.780353e-012, -2.053602e-011,
  2.172643e-014, -8.897365e-015, 2.204596e-011, 3.458929e-011,
  1.147286e-014, -1.411523e-014, 1.997541e-011, 1.804542e-011,
  1.545706e-014, -1.383644e-014, 1.103929e-011, 7.575485e-012,
  1.409382e-014, -1.483454e-014, 1.815812e-011, 1.119613e-011,
  1.570768e-014, -7.939264e-015, 2.938813e-011, 1.299099e-011,
  1.569851e-014, -1.238133e-014, 2.633844e-011, 3.307866e-011,
  2.586231e-014, -6.777544e-015, -8.69737e-012, -2.041628e-011,
  7.916552e-014, -1.900876e-014, -2.415339e-012, 9.604361e-012,
  1.28435e-014, -2.999827e-015, -2.827875e-011, -4.201659e-011,
  2.407412e-014, -1.684545e-014, 7.796671e-012, 1.682111e-011,
  1.740239e-014, -1.091722e-015, 5.156202e-012, -1.638516e-011,
  1.343952e-014, -4.22531e-015, 1.306609e-011, 2.351629e-011,
  9.608732e-015, -4.053112e-015, -2.254696e-011, -3.279556e-011,
  1.699582e-014, 2.75537e-015, 1.286958e-011, 1.143982e-011,
  1.533166e-014, -5.370442e-015, -7.950963e-012, -3.088546e-011,
  1.688753e-014, -1.85648e-015, -9.247647e-012, -3.048265e-012,
  1.264278e-014, -4.814895e-015, 1.164454e-011, -1.369829e-011,
  1.260677e-014, -1.08901e-014, 4.943858e-012, 1.24758e-011,
  1.337382e-014, -1.160605e-014, -2.171771e-011, 2.32861e-012,
  1.600048e-014, -1.305364e-014, 1.109525e-011, 2.358866e-011,
  1.686796e-014, -4.364838e-015, -2.251896e-011, -8.743834e-012,
  1.260657e-014, -1.359168e-014, 2.992351e-011, 2.553518e-011,
  2.489113e-014, -1.832896e-015, -1.061365e-012, -1.253555e-011,
  1.897101e-014, -1.537084e-014, -9.325173e-012, 1.681334e-011,
  3.485144e-014, -1.117644e-014, -1.413581e-011, -2.202804e-012,
  3.17679e-014, -4.88774e-015, -2.2172e-011, -3.436505e-011,
  2.145746e-014, -9.108043e-015, -2.947259e-012, 1.089997e-011,
  1.273392e-014, -8.274606e-015, 1.345447e-011, 2.592539e-011,
  1.014634e-014, -9.52833e-015, -6.459196e-012, -2.332191e-012,
  1.514562e-014, -6.227942e-015, 4.725864e-011, 6.597264e-011,
  1.078465e-014, -5.529359e-015, 1.719885e-011, 4.201312e-011,
  1.014632e-014, -6.088283e-015, 2.297642e-011, 4.098559e-011,
  2.50927e-014, -1.229518e-015, -2.673017e-012, -1.43517e-012,
  2.693481e-014, 1.778837e-015, -6.025246e-013, 1.518604e-011,
  3.576578e-014, -3.638921e-016, -1.164659e-011, -8.571075e-012,
  4.662356e-014, -1.423219e-015, -2.08366e-011, 9.509829e-013,
  5.234938e-014, -1.119108e-015, -3.824288e-012, -3.082942e-012,
  6.50856e-014, -3.530996e-015, -8.22367e-012, 6.438869e-012,
  2.961529e-014, -1.680526e-015, -7.252401e-012, -6.761367e-012,
  2.798911e-014, -5.0432e-016, 1.227327e-011, 2.918499e-011,
  3.403287e-014, -6.149506e-016, -5.859311e-012, -5.18285e-012,
  2.988565e-014, 1.945611e-016, -5.256346e-012, 1.200005e-011,
  3.087528e-014, 6.327378e-016, -1.479019e-011, -2.216257e-011,
  3.272122e-014, 1.118976e-015, 1.877062e-014, 1.03341e-011,
  8.75649e-014, -5.738168e-015, -1.609005e-012, 3.229109e-013,
  8.378884e-014, -4.437628e-015, -2.785277e-013, 1.583497e-011,
  3.280426e-014, 4.316024e-015, 3.050478e-012, 6.453211e-012,
  3.073787e-014, 2.829735e-015, -2.780371e-012, 1.653938e-011,
  3.346455e-014, 3.794634e-015, -7.71984e-012, -1.491447e-012,
  3.553942e-014, 1.748983e-015, -6.456381e-012, 1.168652e-011,
  2.854413e-014, -2.979607e-014, 2.070742e-013, 6.931148e-013,
  4.26948e-014, 5.447562e-014, -1.864691e-012, 1.699907e-011,
  4.978636e-014, -5.824398e-016, 4.906357e-012, 3.194722e-012,
  -3.753104e-014, 1.685073e-014, -5.213582e-012, 1.374144e-011,
  3.414669e-014, 2.60832e-015, 3.170383e-012, 3.657438e-012,
  2.635513e-014, 4.479148e-015, -3.481579e-012, 1.639023e-011,
  3.817911e-014, 3.15874e-015, 1.549162e-012, 4.733744e-012,
  4.0082e-014, 2.922267e-015, -4.3668e-012, 1.883392e-011,
  3.76107e-014, 1.927013e-015, 1.316933e-013, -1.88353e-012,
  3.654428e-014, 3.202926e-015, -3.781971e-012, 1.431728e-011,
  3.950672e-014, 1.529024e-015, 2.631626e-012, 2.734115e-012,
  3.77921e-014, 1.984748e-015, -9.660676e-013, 1.898447e-011,
  4.283262e-014, 4.310074e-015, 1.391891e-012, 2.061831e-012,
  3.849574e-014, 1.571709e-015, 3.016379e-012, 2.485212e-011,
  4.367331e-014, 3.074564e-015, -7.669947e-013, -3.255557e-012,
  4.161674e-014, 1.237938e-015, -1.961868e-011, -3.320097e-012,
  4.336575e-014, 1.844078e-015, -3.253813e-014, -6.373432e-013,
  4.015866e-014, 2.070053e-015, -3.988447e-012, 2.179346e-011,
  4.679003e-014, 7.348683e-015, 5.444394e-012, 7.277314e-012,
  3.935975e-014, -5.246004e-015, -4.818855e-012, 2.037234e-011,
  4.801029e-014, 5.894328e-015, 1.23237e-012, -3.620014e-013,
  4.152038e-014, -1.443709e-015, -2.016252e-012, 2.167362e-011,
  4.570168e-014, 1.911597e-015, -4.048174e-012, -6.145258e-012,
  4.254967e-014, 1.118592e-015, -1.258151e-011, 6.509006e-012,
  4.863756e-014, 4.918302e-016, 1.976127e-013, -2.248987e-012,
  4.799511e-014, -1.040821e-015, 1.79586e-012, 2.424529e-011,
  4.719471e-014, -1.585171e-015, -1.014549e-011, -1.103572e-011,
  4.271707e-014, -1.068563e-015, 1.21477e-011, 3.708837e-011,
  1.440509e-014, 6.287127e-015, 2.429298e-012, 4.373426e-012,
  -6.388927e-014, 1.74674e-014, 1.468337e-011, 3.836011e-011,
  4.940524e-014, -1.55619e-014, -3.921232e-012, 9.26016e-013,
  4.535597e-014, -1.315032e-014, 5.399021e-012, 3.118721e-011,
  5.350595e-014, -1.085148e-014, -4.071215e-012, -2.729629e-012,
  4.790017e-014, -6.437517e-015, 5.162657e-012, 3.128245e-011,
  5.328556e-014, -1.052384e-014, 1.186367e-012, 5.363418e-012,
  5.25097e-014, -9.710665e-015, 1.330886e-012, 3.321207e-011,
  5.894466e-014, -7.147499e-015, 2.422436e-011, 1.796969e-011,
  1.303381e-013, -1.696827e-014, -1.093264e-011, 2.323521e-011,
  6.092175e-014, -6.041528e-015, -8.702779e-012, -9.244942e-012,
  5.900364e-014, -3.560116e-015, 1.086596e-011, 3.857339e-011,
  5.930335e-014, -7.2313e-015, -8.946491e-012, -1.127133e-012,
  5.730767e-014, -7.445597e-015, -7.241611e-012, 1.777467e-011,
  6.158768e-014, -4.249166e-015, -1.818697e-012, -4.292859e-013,
  5.785135e-014, -8.346543e-015, 4.864531e-012, 3.390902e-011,
  6.119169e-014, -5.107092e-015, -4.153124e-012, -6.789477e-011,
  6.539302e-014, -8.306068e-015, 2.970271e-012, 1.267098e-011,
  6.32009e-014, -4.57447e-015, -4.642088e-012, -4.88427e-012,
  6.368024e-014, -6.089483e-015, -1.595843e-011, 1.422015e-011,
  6.338158e-014, -5.062221e-015, 1.116335e-012, 8.589612e-013,
  5.030472e-014, -2.96063e-015, 7.951791e-012, 3.957949e-011,
  6.842303e-014, -1.998379e-015, 1.66527e-012, -2.702699e-012,
  6.679372e-014, -5.214682e-015, 3.245688e-012, 4.32554e-011,
  4.736962e-014, -1.491886e-015, 1.161922e-012, 9.04549e-013,
  9.350612e-014, -1.445433e-014, 8.556445e-012, 5.36378e-011,
  5.792669e-014, -5.8071e-015, 4.17955e-012, 4.951976e-012,
  1.043055e-013, -1.161409e-014, 5.435221e-012, 4.203547e-011,
  7.606994e-014, -8.503729e-015, 2.968922e-012, 6.537726e-013,
  7.453167e-014, -6.279155e-015, 4.063502e-012, 3.909326e-011,
  6.986159e-014, -4.619374e-015, 1.189315e-012, 2.13089e-013,
  7.022028e-014, -3.947415e-015, 1.865752e-012, 4.328587e-011,
  8.190015e-014, -2.7142e-015, -1.970478e-013, -1.534648e-012,
  9.373059e-014, -3.790173e-015, -5.668485e-012, 3.655057e-011,
  1.015845e-013, -3.084722e-015, 4.261158e-012, 1.611344e-012,
  2.01171e-013, -1.802671e-014, -3.451864e-012, 4.111632e-011,
  8.814893e-014, 9.742146e-016, 9.612916e-012, 9.238955e-012,
  9.091245e-014, 1.077308e-015, -6.238038e-012, 4.604334e-011,
  8.613555e-014, 1.303368e-015, 1.201099e-013, -1.510346e-012,
  8.879627e-014, 1.827091e-015, -2.581241e-012, 4.820364e-011,
  9.184189e-014, 3.054317e-015, 2.83398e-013, -7.519719e-014,
  9.199554e-014, 2.798495e-015, -6.906881e-013, 4.955011e-011,
  1.446557e-013, -1.681606e-015, 5.451245e-012, 2.672508e-012,
  3.376099e-014, 1.418162e-014, -2.141067e-012, 5.042267e-011,
  9.289883e-014, 9.569492e-015, 8.586975e-014, -2.641979e-012,
  9.729889e-014, 9.400194e-015, -6.245838e-012, 4.814182e-011,
  9.912234e-014, 1.07917e-014, 3.836399e-012, 4.08929e-012,
  1.023149e-013, 1.154387e-014, -9.804309e-012, 4.703573e-011,
  1.015115e-013, 5.794792e-015, -8.779752e-013, -1.462468e-012,
  1.034425e-013, 8.231527e-015, -5.488604e-012, 5.981143e-011,
  1.37941e-013, -2.090903e-014, 8.552738e-012, 4.436583e-012,
  6.426383e-014, 2.232007e-014, -1.798468e-011, 4.390219e-011,
  1.125051e-013, 1.827581e-014, 4.464205e-012, 3.638818e-012,
  1.079523e-013, 2.508543e-014, 1.073359e-011, 7.490025e-011,
  1.146016e-013, 2.276951e-014, -4.143348e-012, -3.577009e-013,
  1.194467e-013, 2.282882e-014, -4.114763e-012, 6.949935e-011,
  1.182616e-013, 1.779046e-014, 6.297464e-012, 3.787168e-012,
  1.20747e-013, 1.93905e-014, -1.431353e-011, 5.894672e-011,
  1.417396e-013, 1.179135e-014, 2.289201e-012, 1.389108e-012,
  9.018704e-014, 2.085059e-014, -7.514846e-012, 6.45924e-011,
  1.403197e-013, 8.513166e-015, -2.904131e-012, -4.542229e-012,
  1.065546e-013, 2.155505e-014, 1.519771e-012, 7.594722e-011,
  1.366494e-013, 8.368201e-015, 1.703713e-012, 8.431544e-013,
  1.433578e-013, 1.306134e-014, -1.096119e-013, 7.524629e-011,
  1.426226e-013, 6.975025e-015, 5.055162e-012, 3.954497e-012,
  1.459271e-013, 8.006455e-015, -6.042019e-013, 7.605917e-011,
  1.24309e-013, 6.778074e-015, 4.846871e-012, 3.645708e-012,
  1.549072e-013, 4.268982e-015, -5.912375e-012, 7.609597e-011,
  9.905367e-014, 1.087547e-014, -4.101936e-012, -4.805702e-012,
  1.694934e-013, 1.047135e-015, 2.164374e-012, 8.761924e-011,
  1.635992e-013, 1.020154e-016, 2.309005e-012, -6.713716e-014,
  1.678295e-013, 2.547423e-015, -1.509424e-013, 8.604417e-011,
  1.684966e-013, -3.124311e-015, 1.487122e-012, -1.177388e-012,
  1.77584e-013, -2.328653e-015, -2.33912e-012, 8.522733e-011,
  1.774762e-013, -1.052618e-014, -1.565993e-012, -3.84388e-012,
  1.86573e-013, -7.548728e-015, 6.869348e-012, 9.102637e-011,
  1.866678e-013, -1.118837e-014, -9.526639e-013, -3.739474e-012,
  1.923106e-013, -1.14366e-014, 8.183744e-012, 9.56739e-011,
  1.929435e-013, -1.264119e-014, -3.635328e-012, -5.632166e-012,
  2.026141e-013, -1.05561e-014, 6.36679e-012, 9.702895e-011,
  2.024028e-013, -1.233027e-014, -7.257671e-013, -3.817649e-012,
  2.127809e-013, -1.173234e-014, 4.37254e-012, 9.97305e-011,
  2.138565e-013, -1.345236e-014, -1.249952e-012, -8.243027e-012,
  2.238139e-013, -1.300619e-014, 4.7531e-012, 1.067656e-010,
  1.666603e-013, -8.748067e-015, 5.383291e-012, -4.201229e-012,
  2.462386e-013, -1.368991e-014, 8.568556e-012, 1.156479e-010,
  2.331323e-013, -1.574423e-014, -7.480557e-014, -7.548456e-012,
  2.441648e-013, -1.488329e-014, 8.780946e-012, 1.166672e-010,
  2.49495e-013, -1.657184e-014, 5.547397e-012, -8.143541e-012,
  2.567378e-013, -1.210654e-014, -6.906959e-013, 1.184984e-010,
  2.659176e-013, -1.748348e-014, 1.150851e-011, 2.755289e-012,
  2.67051e-013, -1.44605e-014, 1.021737e-012, 1.21438e-010,
  2.625288e-013, -1.034657e-014, 4.231263e-012, -8.959394e-012,
  3.3684e-013, -1.959293e-014, 1.046447e-011, 1.415986e-010,
  2.944432e-013, -1.470677e-014, -5.837771e-013, -1.6622e-011,
  3.148593e-013, -1.293783e-014, 5.178292e-012, 1.474844e-010,
  3.183661e-013, -1.260942e-014, -3.003586e-011, -4.05701e-011,
  3.129883e-013, -1.089212e-014, 7.068832e-013, 1.539824e-010,
  3.364026e-013, -1.686405e-014, 5.402844e-014, -1.859106e-011,
  3.27527e-013, -1.29696e-014, 6.536952e-012, 1.620704e-010,
  3.833544e-013, -2.477734e-014, 1.59555e-012, -1.85579e-011,
  3.578941e-013, -1.802802e-014, 9.927163e-012, 1.729296e-010,
  4.175254e-013, -2.620478e-014, 3.34966e-012, -1.991704e-011,
  3.788552e-013, -1.578318e-014, 6.101066e-012, 1.815703e-010,
  3.993751e-013, -1.225605e-014, 2.442376e-012, -2.425989e-011,
  3.75749e-013, -5.182718e-015, 2.825692e-012, 1.992806e-010,
  4.262407e-013, -9.045346e-015, -7.244078e-013, -2.840465e-011,
  3.920655e-013, 3.8713e-016, 2.370567e-012, 2.109295e-010,
  4.52842e-013, -1.344764e-014, 3.077659e-012, -2.95312e-011,
  4.076401e-013, -1.383383e-015, 8.427192e-012, 2.272741e-010,
  4.778892e-013, -1.877057e-014, 1.014498e-011, -2.267361e-011,
  4.258405e-013, -1.257701e-014, 1.699108e-011, 2.540743e-010,
  5.106035e-013, -2.882804e-014, -9.885774e-012, -5.07001e-011,
  4.466149e-013, -1.982797e-014, 8.522831e-012, 2.572187e-010,
  5.412853e-013, -2.702968e-014, 5.786704e-013, -3.323259e-011,
  4.57334e-013, -2.393278e-014, 5.73867e-012, 2.766384e-010,
  5.690997e-013, -1.902611e-014, 1.301385e-011, -2.41172e-011,
  4.804768e-013, -7.739687e-015, 6.212693e-012, 2.950038e-010,
  6.651268e-013, -1.783041e-014, 7.346017e-012, -3.482513e-011,
  5.29382e-013, -8.98389e-015, 4.538278e-012, 3.33699e-010,
  6.430484e-013, -1.422218e-014, 1.229256e-011, -3.323404e-011,
  5.214664e-013, -1.335229e-014, 8.761455e-012, 3.557813e-010,
  6.791558e-013, -2.563719e-014, 5.675703e-012, -4.765604e-011,
  5.368855e-013, -1.824061e-014, 1.765402e-011, 3.978444e-010,
  7.193272e-013, -2.840873e-014, -3.386734e-012, -5.336569e-011,
  5.620477e-013, -2.199078e-014, 1.621984e-011, 4.314823e-010,
  8.151448e-013, -4.535171e-014, -2.05855e-012, -4.513989e-011,
  5.512969e-013, -1.449819e-014, 1.660621e-011, 4.694428e-010,
  7.995708e-013, -3.403132e-014, 2.127128e-012, -2.919831e-011,
  6.012219e-013, -2.136748e-014, 2.221503e-011, 5.189706e-010,
  8.203248e-013, -4.417705e-014, -5.996809e-014, -2.775289e-011,
  6.372765e-013, -2.954583e-014, 1.781059e-011, 5.513763e-010,
  8.468988e-013, -7.130565e-014, 1.846019e-012, -1.362916e-011,
  6.641725e-013, -5.588807e-014, 1.083891e-011, 5.816093e-010,
  8.256515e-013, -6.240125e-014, -9.826896e-013, -4.577953e-012,
  6.74673e-013, -4.949166e-014, 3.964059e-011, 6.728214e-010,
  8.571123e-013, -5.080404e-014, 1.396915e-011, 4.103629e-011,
  7.280148e-013, -4.235347e-014, 3.710854e-011, 7.420817e-010,
  8.965376e-013, -3.667275e-014, -4.586636e-012, 5.45032e-011,
  7.896727e-013, -2.781992e-014, 2.818455e-011, 8.060467e-010,
  8.956089e-013, -3.079331e-014, 1.545755e-011, 1.002298e-010,
  8.575637e-013, -2.109713e-014, -1.477316e-011, 8.510423e-010,
  8.902054e-013, -3.464025e-014, -2.645564e-012, 1.269684e-010,
  9.356073e-013, -2.861624e-014, 2.247535e-011, 9.608271e-010,
  8.590019e-013, -3.700395e-014, -9.884054e-012, 1.7628e-010,
  1.048939e-012, -4.211822e-014, 3.438772e-011, 1.048118e-009,
  8.142421e-013, -3.795603e-014, 3.145179e-012, 2.613876e-010,
  1.184194e-012, -4.396308e-014, 2.516171e-011, 1.122562e-009,
  7.586131e-013, -2.519489e-014, 7.738865e-012, 3.494316e-010,
  1.362257e-012, -2.686526e-014, 2.707451e-011, 1.223083e-009,
  6.812587e-013, -1.795391e-014, 1.647965e-011, 4.651106e-010,
  1.591006e-012, -1.601446e-014, 1.918149e-011, 1.311035e-009,
  5.86713e-013, -1.639982e-014, 5.984939e-012, 5.680533e-010,
  1.883829e-012, -1.689196e-014, 2.277019e-011, 1.400472e-009,
  4.723151e-013, 6.781097e-015, 5.445253e-012, 7.181016e-010,
  2.269383e-012, 1.940249e-014, 2.148583e-012, 1.484836e-009,
  3.427756e-013, 3.09685e-014, 1.033392e-011, 8.896791e-010,
  2.752825e-012, 5.948168e-014, -1.991074e-011, 1.560095e-009,
  2.274673e-013, 3.190862e-014, 2.241196e-011, 1.096477e-009,
  3.387656e-012, 6.446339e-014, -2.552976e-011, 1.621757e-009,
  4.562239e-014, 3.03471e-014, -1.819621e-011, 1.276089e-009,
  4.192651e-012, 4.183302e-014, -1.480395e-011, 1.655735e-009,
  -8.817205e-014, 3.114726e-014, 1.961193e-011, 1.559716e-009,
  5.201057e-012, 3.241505e-014, 1.011053e-011, 1.671701e-009,
  -1.637128e-013, 2.542372e-014, 1.770349e-011, 1.858063e-009,
  6.404238e-012, 3.093367e-014, -2.892194e-011, 1.638716e-009,
  -2.284048e-013, 2.261728e-014, 2.709541e-011, 2.19526e-009,
  8.14305e-012, -1.928013e-015, -9.345947e-012, 1.584631e-009,
  -1.610064e-013, -3.736463e-014, 3.135223e-011, 2.545163e-009,
  1.021503e-011, -1.181259e-013, 1.094597e-011, 1.432427e-009,
  7.314735e-014, -1.359812e-013, 5.298362e-011, 2.927272e-009,
  1.282105e-011, -3.03005e-013, 4.896085e-011, 1.187254e-009,
  5.844762e-013, -1.524913e-013, 6.629995e-011, 3.330074e-009,
  1.607444e-011, -3.24324e-013, 4.578261e-011, 8.459253e-010,
  1.508621e-012, -1.938554e-013, 6.402812e-011, 3.729582e-009,
  2.016537e-011, -3.675032e-013, 4.560911e-011, 3.641351e-010,
  3.048233e-012, -3.402048e-013, 8.563263e-011, 4.123291e-009,
  2.524123e-011, -5.55203e-013, 6.791354e-011, -3.144946e-010,
  5.462377e-012, -6.465682e-013, 1.236354e-010, 4.450028e-009,
  3.16478e-011, -9.245687e-013, 1.132847e-010, -1.249595e-009,
  9.12752e-012, -1.026785e-012, 1.719244e-010, 4.665448e-009,
  3.960138e-011, -1.295375e-012, 1.453635e-010, -2.496445e-009,
  1.456957e-011, -1.595064e-012, 2.170009e-010, 4.670388e-009,
  4.965338e-011, -1.749741e-012, 1.763772e-010, -4.158353e-009,
  2.256297e-011, -2.228917e-012, 2.596029e-010, 4.365091e-009,
  6.228626e-011, -2.110779e-012, 2.198642e-010, -6.298205e-009,
  3.437182e-011, -3.657546e-012, 3.356673e-010, 3.55771e-009,
  7.798114e-011, -2.995778e-012, 2.828017e-010, -9.102834e-009,
  5.150541e-011, -5.600775e-012, 4.433811e-010, 2.016016e-009,
  9.760712e-011, -4.044204e-012, 3.62351e-010, -1.266055e-008,
  7.689058e-011, -7.07592e-012, 4.220283e-010, -6.690204e-010,
  1.206234e-010, -4.565048e-012, 3.274693e-010, -1.72576e-008,
  1.149316e-010, -9.58934e-012, 4.291796e-010, -5.152045e-009,
  1.520169e-010, -4.788706e-012, 3.692777e-010, -2.315507e-008,
  1.706724e-010, -1.425319e-011, 5.512042e-010, -1.244443e-008,
  1.927062e-010, -5.929748e-012, 5.201861e-010, -3.087705e-008,
  2.560476e-010, -1.88437e-011, 6.217345e-010, -2.428576e-008,
  2.448575e-010, -6.348006e-012, 6.357641e-010, -4.099358e-008,
  3.88956e-010, -2.408113e-011, 6.272504e-010, -4.329782e-008,
  3.119234e-010, -6.145669e-012, 7.310071e-010, -5.408619e-008,
  6.073247e-010, -3.035749e-011, 7.581518e-010, -7.50706e-008,
  4.028372e-010, -5.241045e-012, 9.215561e-010, -7.177049e-008,
  9.79958e-010, -3.767105e-011, 1.404683e-009, -1.293955e-007,
  5.271209e-010, -2.493332e-012, 1.516013e-009, -9.561396e-008,
  1.655852e-009, -6.081486e-011, 4.281611e-009, -2.30581e-007,
  6.985429e-010, 2.500478e-012, 3.131059e-009, -1.296381e-007,
  2.868374e-009, -1.174301e-010, 1.217311e-008, -4.389223e-007,
  9.32157e-010, 8.964029e-012, 6.177378e-009, -1.7992e-007,
  4.019476e-009, -2.766053e-010, 3.615083e-008, -9.364401e-007,
  1.154855e-009, 1.941456e-011, 1.181124e-008, -2.590654e-007,
  -1.141954e-009, -5.830758e-010, 1.034899e-007, -2.114697e-006,
  1.077891e-009, 3.210944e-011, 2.178415e-008, -3.74111e-007,
  -1.093877e-008, -6.13068e-010, 1.64042e-007, -3.504447e-006,
  1.1157e-009, 4.448318e-011, 2.642699e-008, -4.638751e-007,
  -1.294965e-008, -6.053067e-010, 1.634299e-007, -3.917238e-006,
  1.179996e-009, 2.596718e-011, 2.24029e-008, -4.825213e-007,
  -9.945849e-009, -1.023497e-009, 1.106896e-007, -3.295809e-006,
  1.305396e-009, -1.863617e-011, 1.545992e-008, -4.192882e-007,
  2.927437e-010, -1.10019e-009, 4.603903e-008, -1.876783e-006,
  1.408777e-009, -1.595498e-011, 9.928644e-009, -3.077436e-007,
  4.082721e-009, -4.439517e-010, 1.636747e-008, -8.318423e-007,
  1.124882e-009, 1.359776e-012, 6.105814e-009, -2.226464e-007,
  2.721446e-009, -9.459733e-011, 5.460542e-009, -3.99705e-007,
  8.604651e-010, 5.049023e-012, 2.907057e-009, -1.625538e-007,
  1.565522e-009, -1.710254e-011, 1.40087e-009, -2.149655e-007,
  6.510866e-010, 9.266207e-013, 1.110287e-009, -1.205989e-007,
  9.314307e-010, -2.049292e-011, 5.754422e-010, -1.226423e-007,
  4.955562e-010, -3.716611e-012, 6.449191e-010, -9.051404e-008,
  5.831727e-010, -2.613432e-011, 5.338385e-010, -7.235762e-008,
  3.838243e-010, -7.693682e-012, 6.414966e-010, -6.885966e-008,
  3.789742e-010, -2.981517e-011, 9.097254e-010, -4.297464e-008,
  3.008131e-010, -9.802219e-012, 8.835874e-010, -5.287008e-008,
  2.517123e-010, -2.392371e-011, 9.768878e-010, -2.501883e-008,
  2.37679e-010, -8.85358e-012, 9.462544e-010, -4.057172e-008,
  1.700963e-010, -1.519985e-011, 8.465098e-010, -1.368981e-008,
  1.896534e-010, -6.539969e-012, 8.05149e-010, -3.123625e-008,
  1.163099e-010, -7.941895e-012, 6.438121e-010, -6.452797e-009,
  1.517795e-010, -3.979274e-012, 6.170835e-010, -2.389299e-008,
  7.947048e-011, -6.31317e-012, 5.835211e-010, -1.940922e-009,
  1.219618e-010, -3.99618e-012, 6.360298e-010, -1.816406e-008,
  5.386447e-011, -4.773373e-012, 5.969336e-010, 9.065476e-010,
  9.910819e-011, -3.331726e-012, 6.332624e-010, -1.372186e-008,
  3.652737e-011, -4.045882e-012, 5.165304e-010, 2.529112e-009,
  7.995297e-011, -3.11945e-012, 6.510033e-010, -1.02101e-008,
  2.454079e-011, -2.856234e-012, 4.249443e-010, 3.475321e-009,
  6.45351e-011, -2.29039e-012, 5.669243e-010, -7.433171e-009,
  1.613602e-011, -1.442258e-012, 2.441274e-010, 3.954699e-009,
  5.204634e-011, -1.059472e-012, 3.963364e-010, -5.23171e-009,
  1.039667e-011, -1.69016e-013, 7.653575e-011, 4.105122e-009,
  4.194085e-011, 1.244005e-013, 1.836882e-010, -3.530209e-009,
  6.446892e-012, -1.108171e-013, 7.152232e-011, 4.056863e-009,
  3.377039e-011, 3.39007e-014, 1.563443e-010, -2.197869e-009,
  3.773406e-012, -3.142567e-013, 1.004687e-010, 3.852217e-009,
  2.718147e-011, -2.506782e-013, 2.25025e-010, -1.088321e-009,
  1.989255e-012, -2.239603e-013, 9.066705e-011, 3.593744e-009,
  2.189636e-011, -1.470098e-013, 1.290783e-010, -3.72181e-010,
  8.680401e-013, -1.035227e-013, 6.082117e-011, 3.268845e-009,
  1.768371e-011, 4.271804e-014, 1.016823e-010, 2.597576e-010,
  1.837711e-013, -7.4704e-014, 9.725655e-012, 2.911036e-009,
  1.426255e-011, 7.523165e-014, 6.657042e-011, 6.602566e-010,
  -1.608006e-013, -8.845153e-014, 5.334026e-011, 2.634289e-009,
  1.158597e-011, -1.480186e-014, 8.432842e-011, 9.864785e-010,
  -3.465284e-013, -5.280665e-014, 1.846802e-011, 2.283222e-009,
  9.33136e-012, -2.415371e-015, 8.089526e-011, 1.201602e-009,
  -3.837902e-013, -3.274486e-014, -4.594689e-011, 1.904509e-009,
  7.588402e-012, 5.694232e-014, 4.225558e-011, 1.327363e-009,
  -3.336292e-013, -1.523853e-014, -2.174275e-011, 1.669271e-009,
  6.145731e-012, 7.976084e-014, -8.660169e-012, 1.368737e-009,
  -2.351848e-013, -4.557952e-015, -1.31554e-012, 1.467545e-009,
  5.011383e-012, 5.107739e-014, 1.13659e-011, 1.425992e-009,
  -1.259686e-013, -2.826303e-014, 2.565161e-012, 1.239124e-009,
  4.10717e-012, 2.341187e-014, 7.429463e-012, 1.406545e-009,
  9.688755e-015, -3.303606e-014, 6.940367e-012, 1.041865e-009,
  3.374014e-012, -5.858667e-016, -1.955672e-012, 1.37632e-009,
  1.430252e-013, -3.180445e-014, 7.710066e-013, 8.687571e-010,
  2.790615e-012, -2.207013e-014, 2.369885e-011, 1.355329e-009,
  2.572928e-013, -3.862676e-014, 1.808754e-011, 7.314076e-010,
  2.325491e-012, 3.193174e-015, -7.982916e-012, 1.273907e-009,
  3.693619e-013, 2.324949e-014, -1.948024e-012, 5.928516e-010,
  1.95576e-012, 6.354114e-014, -3.118776e-011, 1.238281e-009,
  4.617082e-013, 3.636309e-014, 1.339287e-012, 4.83141e-010,
  1.660541e-012, 9.045169e-014, -4.877797e-011, 1.170682e-009,
  5.406882e-013, 2.577611e-014, -1.280727e-011, 3.740501e-010,
  1.421155e-012, 8.074113e-014, -4.950202e-011, 1.090259e-009,
  6.051948e-013, 1.768425e-014, -2.1221e-011, 2.819256e-010,
  1.240092e-012, 4.026568e-014, -2.878331e-011, 1.024375e-009,
  6.570367e-013, -2.957379e-014, 3.402453e-012, 2.445549e-010,
  1.082122e-012, -3.261219e-014, 3.2372e-011, 9.723696e-010,
  6.907362e-013, -5.807905e-014, 3.708327e-012, 1.780285e-010,
  9.673146e-013, -7.552012e-014, 2.975292e-011, 8.625528e-010,
  7.137523e-013, -7.477845e-014, -2.355709e-011, 9.98413e-011,
  8.761006e-013, -5.558353e-014, 3.693001e-011, 7.9709e-010,
  7.290636e-013, 3.90697e-015, -2.209095e-012, 9.245568e-011,
  7.90923e-013, -5.925155e-014, 4.069604e-011, 7.916552e-010,
  7.046386e-013, 2.282432e-014, -2.890459e-011, 1.452427e-011,
  7.984485e-013, -3.275287e-016, 2.932772e-011, 7.506646e-010,
  7.21076e-013, -4.743128e-014, -5.376873e-011, -3.912904e-011,
  6.921502e-013, 5.162741e-015, -4.598742e-011, 5.642379e-010,
  7.223257e-013, -7.421239e-015, -2.689835e-011, -1.251607e-011,
  6.489987e-013, -9.78595e-015, 1.078411e-012, 5.950436e-010,
  7.142886e-013, -1.057054e-015, -1.895276e-011, -2.335189e-011,
  6.139517e-013, -2.062454e-014, 1.539629e-011, 5.750657e-010,
  7.350671e-013, 5.138328e-015, -1.196671e-011, -2.321612e-011,
  6.35831e-013, -2.805256e-014, 4.57412e-011, 5.6912e-010,
  6.869708e-013, -3.526928e-014, 2.213798e-011, 6.91642e-012,
  5.720363e-013, -2.861744e-014, 3.868121e-011, 4.960032e-010,
  6.588191e-013, -4.598392e-014, 9.89432e-012, -1.710104e-012,
  5.417914e-013, -5.334068e-014, 3.714237e-011, 4.511749e-010,
  6.312254e-013, -6.159269e-014, -1.512732e-011, -4.472799e-011,
  5.251403e-013, -5.387214e-014, 3.603257e-011, 4.046311e-010,
  6.256275e-013, -5.041933e-014, 6.585894e-013, -4.323946e-011,
  4.645854e-013, -4.367148e-014, 3.652353e-011, 3.795406e-010,
  5.859698e-013, -6.210072e-014, -1.928022e-011, -6.05118e-011,
  4.598275e-013, -5.477119e-014, 4.581774e-011, 3.616449e-010,
  5.538422e-013, -8.737884e-014, 1.769062e-011, -1.004203e-011,
  4.777405e-013, -7.579977e-014, 5.993698e-011, 3.237903e-010,
  5.227397e-013, -7.840047e-014, 1.057587e-011, -1.947571e-011,
  4.520084e-013, -8.001605e-014, 7.00982e-011, 3.208173e-010,
  4.959965e-013, -4.714844e-014, -2.590717e-011, -8.341153e-011,
  4.44531e-013, -1.504739e-014, 2.006321e-011, 2.62319e-010,
  4.853679e-013, -2.405362e-014, -1.782172e-011, -5.127894e-011,
  4.298723e-013, -2.915279e-014, 4.023522e-011, 2.87204e-010,
  4.584657e-013, -2.325006e-014, -4.682069e-011, -8.027159e-011,
  4.025213e-013, -2.51465e-014, 5.119424e-011, 2.969425e-010,
  4.312056e-013, -5.25156e-015, 3.782934e-012, -1.558468e-011,
  3.833102e-013, -5.314443e-014, 4.50049e-011, 2.69667e-010,
  4.105067e-013, -3.774822e-014, 9.038853e-012, -2.346017e-011,
  3.766658e-013, -3.056676e-014, -9.02148e-012, 1.657893e-010,
  4.441306e-013, -7.595118e-014, -2.792499e-011, -6.481322e-011,
  3.355147e-013, -4.118021e-014, 3.988612e-011, 2.195845e-010,
  3.721005e-013, -5.080521e-014, -2.427121e-012, -2.520162e-011,
  3.503736e-013, -4.893574e-014, 4.507484e-011, 1.961784e-010,
  3.553686e-013, -7.410284e-014, -1.344348e-011, -3.041372e-011,
  3.282065e-013, -1.007651e-013, 4.819566e-011, 1.870848e-010,
  3.288784e-013, -7.73578e-014, -1.286052e-011, -6.043228e-011,
  3.24661e-013, -4.326359e-014, 2.582058e-011, 1.540026e-010,
  3.171953e-013, -1.000079e-013, 6.904237e-012, 4.585804e-012,
  2.323747e-013, -9.04466e-014, 4.242457e-011, 1.436813e-010,
  2.941482e-013, -8.829694e-014, -2.145855e-011, -3.147337e-011,
  2.854938e-013, -1.010895e-013, 3.02583e-011, 1.24428e-010,
  2.770553e-013, -9.372769e-014, -1.377455e-011, -2.362498e-011,
  2.75648e-013, -1.018687e-013, 3.053011e-011, 1.120073e-010,
  2.628332e-013, -8.428916e-014, -1.266298e-012, -1.177066e-011,
  2.649672e-013, -8.803735e-014, 1.759113e-011, 9.243294e-011,
  2.048157e-013, -4.31102e-014, -1.855752e-011, -1.782493e-011,
  2.860966e-013, -5.942188e-014, 3.280616e-011, 1.348388e-010,
  2.226752e-013, -3.737171e-014, -1.932013e-011, -4.04464e-011,
  2.584805e-013, -4.16047e-014, 8.894528e-013, 9.899868e-011,
  2.2654e-013, -3.544495e-014, -1.670914e-011, -4.023506e-011,
  2.407874e-013, -2.764826e-014, 8.813966e-012, 1.057271e-010,
  2.150483e-013, -3.111858e-014, -2.457461e-012, -1.967327e-011,
  2.296681e-013, -2.850082e-014, 1.56932e-011, 1.102479e-010,
  2.022133e-013, -4.19453e-014, 2.246213e-012, 6.265408e-012,
  2.154993e-013, -3.976213e-014, 1.950914e-011, 9.812599e-011,
  1.935515e-013, -1.467858e-014, 6.992245e-012, 1.742313e-012,
  2.038886e-013, -3.865457e-014, 2.701563e-011, 1.19522e-010,
  1.889372e-013, -3.412794e-014, -9.817883e-012, -2.679229e-011,
  1.997685e-013, -3.518163e-014, 1.14364e-011, 9.475627e-011,
  1.781098e-013, -4.424669e-014, 5.507522e-013, 3.539543e-012,
  1.875383e-013, -4.565561e-014, 2.073388e-011, 8.989896e-011,
  1.498898e-013, -7.744848e-014, -8.006823e-013, 1.988967e-011,
  1.769545e-013, -5.628515e-014, 4.984855e-012, 4.940311e-011,
  1.077742e-013, -1.228109e-014, -4.465763e-012, 1.628908e-011,
  1.597495e-013, -6.754459e-014, 3.15557e-012, 7.462945e-011,
  1.57125e-013, 1.065086e-014, -3.772904e-012, -3.38252e-013,
  1.623616e-013, -3.809569e-014, 4.521507e-011, 1.422173e-010,
  1.485066e-013, -5.702927e-015, 4.861135e-011, 6.783083e-011,
  1.567496e-013, -2.712545e-014, 6.362722e-011, 1.471993e-010,
  1.408305e-013, -2.019035e-014, 4.519218e-011, 4.052609e-011,
  1.495087e-013, -2.763507e-014, -2.691765e-011, 7.539667e-012,
  8.97405e-014, 1.299866e-014, -2.499851e-011, -4.651034e-011,
  2.036176e-013, 9.185617e-015, -1.236503e-011, 3.859318e-011,
  1.318613e-013, -3.064591e-015, -3.518149e-011, -7.311805e-011,
  1.431416e-013, 1.856797e-014, -3.816254e-011, 1.862278e-012,
  1.301216e-013, -3.413736e-014, -4.864075e-011, -6.147682e-011,
  1.306005e-013, -4.205991e-014, -1.921613e-011, 3.523588e-011,
  1.186483e-013, -3.688462e-014, -2.155469e-011, -2.358187e-011,
  1.346351e-013, -1.205607e-014, 4.033377e-011, 9.767407e-011,
  1.702283e-013, -6.478952e-014, -6.906899e-011, -7.383447e-011,
  1.505873e-013, -9.555365e-015, -3.963362e-011, -2.602683e-011,
  1.287671e-013, -6.003316e-014, 8.678509e-011, 1.252646e-010,
  1.13175e-013, -4.493112e-014, 4.16013e-011, 4.673644e-011,
  9.320457e-014, -4.361418e-014, 2.90295e-011, 1.014758e-011,
  1.169447e-013, -2.674082e-014, -1.058695e-010, -1.123025e-010,
  1.003326e-013, -6.980364e-014, 2.727026e-011, 4.677353e-011,
  1.054782e-013, -5.600657e-014, -4.381938e-011, -2.728539e-011,
  1.351651e-013, -7.758546e-014, -2.837405e-011, -7.296068e-011,
  1.173937e-013, -1.094304e-014, -4.763006e-013, -6.411081e-012,
  1.08991e-013, -6.060709e-014, 3.948415e-011, 5.241396e-011,
  1.044757e-013, -3.940287e-014, 3.143665e-011, 4.008894e-011,
  8.489391e-014, -3.402802e-014, -5.442461e-011, -6.684885e-011,
  1.048657e-013, -1.037896e-014, 3.849797e-011, 8.595166e-011,
  8.786733e-014, -3.280518e-014, 7.469017e-012, -2.829349e-011,
  9.332267e-014, -3.355136e-014, 1.21801e-011, 4.795515e-011,
  1.033114e-013, -2.691933e-014, 2.311857e-011, 2.139954e-011,
  7.459978e-014, -2.84119e-014, 1.718085e-011, 4.499776e-011,
  1.197071e-013, -2.490559e-014, 3.790048e-011, 5.855592e-011,
  4.479741e-014, -4.795828e-014, 8.395456e-012, 1.831779e-011,
  8.719857e-014, -4.795137e-014, -1.566056e-011, -1.420907e-011,
  9.101864e-014, -3.281959e-014, 6.174578e-013, 3.496349e-011,
  8.419759e-014, -1.72187e-014, 4.942955e-011, 4.859159e-011,
  8.443812e-014, -3.059604e-014, 2.220856e-011, 4.991374e-011,
  7.82316e-014, -2.541255e-014, -1.699942e-012, 2.808126e-012,
  7.861135e-014, -3.282801e-014, -1.572897e-011, 1.915601e-011,
  1.859117e-014, -1.153953e-014, -2.463465e-011, -1.158488e-011,
  2.905194e-014, -3.009541e-014, 8.292613e-012, 4.126884e-011,
  6.90037e-014, -2.47702e-014, -5.739163e-012, -6.388833e-013,
  8.047335e-014, -3.690778e-014, 2.682438e-011, 4.89814e-011,
  6.935538e-014, -2.025673e-014, 5.497853e-013, -1.875209e-012,
  7.78861e-014, -2.264068e-014, 2.021153e-011, 4.527387e-011,
  6.578931e-014, -1.736044e-014, 5.492915e-013, 4.012435e-013,
  7.106093e-014, -2.504612e-014, 2.631241e-011, 5.4955e-011,
  6.651427e-014, -2.419841e-014, 4.319435e-012, 4.487994e-013,
  7.259217e-014, -2.546223e-014, 7.566743e-012, 3.090381e-011,
  6.420586e-014, -3.382897e-014, -3.401978e-012, -5.761524e-012,
  6.875209e-014, -2.669064e-014, 8.546086e-012, 2.150199e-011,
  6.443666e-014, -2.980091e-014, -3.471096e-012, -1.091545e-011,
  6.906178e-014, -2.718232e-014, 1.302228e-011, 3.257969e-011,
  5.082422e-014, -3.037226e-014, -1.42637e-011, -1.874267e-011,
  8.715037e-014, -2.789716e-014, 2.444181e-011, 4.095394e-011,
  1.004641e-014, -1.317808e-014, 5.080207e-012, 1.000892e-011,
  7.218485e-014, -3.335417e-014, 2.293136e-011, 3.882857e-011,
  3.616463e-014, -1.639425e-014, -1.905292e-011, -2.277632e-011,
  6.831565e-014, -3.851839e-014, 3.123958e-011, 6.186861e-011,
  1.063658e-014, -1.422046e-014, 1.104062e-012, -7.18796e-012,
  9.334194e-014, -1.049551e-014, 1.900103e-011, 4.207558e-011,
  4.344517e-014, -1.961686e-014, -1.302799e-011, -1.485684e-011,
  7.018719e-014, -2.723832e-014, 1.959128e-011, 3.261183e-011,
  6.904367e-014, -1.96767e-014, -7.469923e-012, -1.324296e-011,
  7.57365e-014, -2.777659e-014, 2.868726e-011, 4.065103e-011,
  9.408602e-014, -2.781622e-014, 9.564569e-012, 8.744326e-012,
  8.690549e-014, -2.816443e-014, 4.510607e-011, 5.64433e-011,
  4.933602e-014, -3.441141e-014, -7.431084e-012, -8.528118e-012,
  5.615713e-014, -2.066713e-014, 2.283879e-011, 2.462532e-011,
  4.721004e-014, -2.595781e-014, 8.461951e-012, 1.986151e-012,
  5.206422e-014, -2.990229e-014, -3.511052e-011, -3.289916e-011,
  4.581398e-014, -2.611945e-014, -3.366655e-011, -3.563808e-011,
  4.858246e-014, -3.057696e-014, 1.454429e-011, 3.554465e-011,
  5.325127e-014, -9.309469e-015, 4.470117e-011, 4.632727e-011,
  4.418655e-014, -1.469246e-014, 8.567717e-011, 1.109819e-010,
  4.762778e-014, -7.885013e-015, -3.332807e-012, -2.086275e-012,
  4.218077e-014, -1.48e-014, 2.342404e-011, 3.258946e-011,
  4.594188e-014, -1.467696e-014, 1.240231e-012, -5.385256e-012,
  5.184783e-014, -1.380215e-014, 3.508211e-012, 3.85728e-012,
  4.655715e-014, 1.305174e-014, -2.557993e-011, -4.393223e-011,
  5.664723e-014, 3.040738e-017, 2.726134e-011, 5.692288e-011,
  1.14732e-013, -8.673451e-015, 1.436615e-011, 5.526576e-012,
  2.067987e-014, 1.962548e-014, 3.085299e-011, 5.685654e-011,
  4.315153e-014, -9.552509e-015, 3.699446e-011, 1.269043e-011,
  5.08337e-014, -5.28477e-015, 2.771792e-011, 4.055496e-011,
  4.786698e-014, 6.405713e-015, 5.024405e-012, 7.195138e-015,
  2.479797e-014, -1.840838e-014, 2.86457e-011, 4.285753e-011,
  5.117503e-014, -4.702646e-015, -5.747175e-011, -5.955753e-011,
  5.80185e-014, -4.560526e-014, 2.429817e-011, 5.740891e-011,
  4.117643e-014, 8.324716e-016, -5.216307e-012, 1.286285e-011,
  -1.436438e-014, -1.806003e-014, -2.417548e-011, 1.096731e-012,
  4.535423e-014, -1.206623e-014, -2.304397e-011, -4.666988e-011,
  1.801473e-014, -1.394923e-014, 2.394769e-011, 6.807319e-011,
  4.40543e-014, -2.266935e-014, -7.214541e-011, -7.611056e-011,
  3.872123e-014, -2.400163e-015, 4.47468e-011, 5.633658e-011,
  4.59871e-014, 3.583914e-014, 2.0108e-011, 2.338798e-011,
  4.504971e-014, -2.074172e-014, 1.184918e-010, 1.705415e-010,
  3.476157e-014, -1.803865e-014, -1.240782e-013, -9.416089e-012,
  3.419313e-014, -2.434785e-014, 7.955626e-011, 1.203094e-010,
  5.124787e-014, -3.040169e-014, 2.875696e-011, 2.39748e-011,
  4.333074e-014, -9.655916e-015, -2.797449e-011, -1.313639e-011,
  3.419817e-014, -1.085318e-014, -2.140621e-011, -2.647584e-011,
  3.050741e-014, -2.509918e-015, 3.336927e-011, 4.514355e-011,
  3.32087e-014, -2.414309e-014, -4.310175e-012, -1.922375e-011,
  2.661967e-014, 2.459823e-015, -2.897854e-012, 5.48461e-012,
  2.144904e-014, -1.505246e-014, -1.402117e-011, -3.963231e-011,
  2.901341e-014, 2.587244e-015, -2.06631e-011, -1.255037e-011,
  -3.365615e-014, -1.298609e-014, -1.444618e-011, -2.348264e-011,
  1.052341e-014, -1.530012e-014, -2.204114e-012, -5.117646e-012,
  3.351017e-014, -2.4167e-014, -4.658781e-012, -1.158992e-011,
  2.653133e-014, -2.098341e-014, 4.199711e-011, 5.54485e-011,
  2.496174e-014, -1.445812e-014, -3.91447e-011, -5.47365e-011,
  3.316666e-014, -1.489727e-014, -2.310465e-011, -1.754087e-011,
  2.870028e-014, -6.926414e-015, -6.178003e-012, -1.037693e-011,
  3.34137e-014, -1.289577e-014, -1.69021e-011, -1.116633e-011,
  4.350637e-014, -1.834874e-014, 7.43672e-012, 6.527026e-012,
  1.034387e-013, -2.583255e-014, 8.278306e-012, 5.353764e-012,
  2.441443e-014, -8.576389e-015, 3.713123e-011, 3.079419e-011,
  2.555551e-014, 6.77745e-015, -1.066473e-011, -9.04271e-012,
  2.495604e-014, -1.49512e-014, -2.101184e-011, -3.24791e-011,
  2.866426e-014, -7.417692e-015, 2.518865e-012, 1.270661e-011,
  1.903289e-014, -2.333079e-014, -4.228185e-012, 2.884229e-011,
  1.699499e-014, -5.098857e-014, 7.590761e-012, 1.572322e-011,
  2.646467e-014, -1.18904e-014, -5.498115e-012, 5.575851e-012,
  1.680422e-014, -2.98638e-014, 4.400642e-011, 5.395275e-011,
  3.101433e-014, -3.551932e-015, -5.257714e-011, -5.847789e-011,
  1.991785e-014, -1.836433e-014, -2.909606e-011, -2.528996e-011,
  1.742248e-014, -4.675556e-014, 7.181285e-011, 1.01571e-010,
  1.8904e-014, -1.205754e-015, 2.192234e-012, -1.188491e-011,
  2.397878e-014, -2.184144e-014, -5.862126e-012, -1.321134e-011,
  2.726792e-014, -1.285322e-014, 1.658502e-011, 1.059422e-011,
  2.000214e-014, -4.382029e-014, 5.42941e-012, 2.838275e-011,
  2.234705e-014, -4.019854e-014, 7.612379e-012, -2.840931e-014,
  3.611881e-014, -3.805557e-015, -2.632499e-012, 1.869129e-011,
  2.041295e-014, -1.903346e-014, 5.949977e-011, 8.588951e-011,
  2.417645e-014, -1.23939e-014, -3.584841e-012, -2.775212e-011,
  2.467894e-014, -3.607418e-015, 2.758218e-011, 3.22407e-011,
  2.442827e-014, -6.69048e-015, -9.017557e-012, -1.353844e-011,
  2.492345e-014, -6.753925e-015, 6.465206e-012, 8.769623e-012,
  3.332647e-014, 3.755002e-015, -4.805745e-011, -5.225347e-011,
  2.910597e-014, -8.802372e-015, -1.211246e-011, 1.391497e-012,
  4.359816e-014, -3.684094e-014, -1.692527e-011, -1.95129e-012,
  6.07696e-014, -2.917066e-014, -2.003397e-011, -4.828995e-011,
  2.198026e-014, -2.592347e-014, 1.071417e-011, -5.108415e-012,
  2.867061e-014, -1.367531e-016, -4.250745e-011, -6.29376e-011,
  2.415971e-014, -4.73248e-015, -1.054089e-011, -1.382233e-011,
  2.313694e-014, -1.739104e-014, 5.535502e-011, 7.069793e-011,
  1.746927e-014, -1.217273e-014, 4.967379e-012, 1.406567e-011,
  1.903957e-014, -2.027156e-015, 1.350956e-011, 5.38193e-011,
  4.956576e-014, 3.90888e-015, 3.826675e-012, 8.021407e-012,
  -4.364328e-014, -1.109446e-014, 2.391982e-011, 4.522439e-011,
  1.659671e-014, -2.058556e-015, 2.036168e-011, 1.376058e-011,
  2.434182e-014, -1.90426e-015, -6.168445e-012, -3.882949e-012,
  2.299623e-014, 1.377247e-014, -1.482563e-011, -1.427071e-011,
  1.827404e-014, -3.227195e-014, 1.280392e-011, 3.932852e-011,
  2.030417e-014, -8.118856e-015, -1.25685e-011, -1.622939e-011,
  1.160332e-014, -1.582826e-014, 3.828044e-011, 5.243308e-011,
  1.790057e-014, -1.092477e-014, 4.601826e-011, 8.76471e-011,
  6.402934e-015, -5.62816e-014, 3.678524e-011, 5.150456e-011,
  1.715779e-014, -5.834262e-015, 1.331267e-011, 1.540639e-011,
  2.268436e-014, -6.903227e-015, 2.780039e-011, 3.567677e-011,
  7.563319e-015, -2.029049e-014, -5.361176e-012, -2.860471e-011,
  2.645619e-014, 1.723623e-014, -2.7857e-011, -2.482057e-011,
  6.134318e-015, -7.113167e-016, -2.070587e-011, -4.895069e-011,
  2.812733e-014, 3.14474e-015, -3.772707e-011, -5.462627e-011,
  -2.837068e-014, -2.134474e-014, -2.666472e-011, -2.051877e-011,
  -2.783143e-014, -1.725507e-014, 3.717503e-011, 2.755194e-011,
  6.633213e-015, -8.229638e-015, -5.53188e-012, -1.137806e-011,
  5.150814e-015, -3.730564e-014, 3.155601e-011, 5.744753e-011,
  1.50972e-014, -3.652955e-014, -3.223176e-011, -4.289228e-011,
  2.079278e-014, -2.845971e-014, -5.278017e-011, -4.309359e-011,
  1.892013e-014, -3.30325e-014, -1.2815e-011, -5.378336e-011,
  5.46627e-015, -2.175309e-014, 6.52127e-011, 7.167944e-011,
  -1.843022e-015, 1.436828e-014, 2.650453e-011, -1.778561e-013,
  3.039995e-014, 2.829115e-014, -8.982729e-012, 6.707567e-012,
  -2.767081e-014, 5.21808e-015, -5.76384e-011, -6.588552e-011,
  3.847083e-014, -1.079774e-014, 3.940882e-011, 7.619263e-011,
  3.314897e-014, -1.704535e-014, 4.502976e-011, 5.831039e-011,
  1.190794e-014, 4.239505e-015, 1.690686e-011, -1.256496e-011,
  2.590567e-014, 1.135398e-016, -2.612432e-011, -3.238907e-011,
  2.405001e-014, -6.644522e-015, 5.391642e-012, 9.564739e-012,
  8.607087e-015, -3.449511e-014, 6.362853e-013, -1.301411e-012,
  8.689044e-015, -1.35698e-014, 2.195118e-012, 2.016877e-011,
  9.954389e-015, -4.671156e-015, 2.5687e-011, 5.897829e-011,
  4.731625e-016, -2.927161e-014, -1.327586e-011, -1.891262e-012,
  1.932495e-014, 1.296447e-015, 2.490173e-011, 4.841089e-011,
  1.031229e-014, -8.150314e-016, 2.566068e-011, 3.151304e-011,
  1.853821e-014, -2.945293e-016, 3.937637e-011, 5.230076e-011,
  1.612658e-014, 7.573403e-015, 2.857895e-011, 3.672415e-011,
  1.574324e-014, -2.461598e-014, -3.869874e-012, -3.380403e-011,
  1.33359e-014, -1.190348e-014, -2.625332e-011, -2.129885e-011,
  1.059141e-014, -1.944149e-014, -2.604755e-011, -4.272255e-011,
  9.113413e-014, -1.73028e-014, 6.917949e-011, 8.075037e-011,
  1.368725e-014, 8.162842e-015, -1.709438e-012, -1.269661e-011,
  2.044456e-014, 2.302028e-014, 6.522374e-011, 1.06834e-010,
  3.389138e-015, -1.416741e-014, -1.243357e-013, -3.52034e-012,
  1.073471e-014, -9.598243e-015, 1.437105e-011, 1.191966e-011,
  1.149905e-014, -3.043737e-014, 2.046847e-011, 2.856078e-011,
  6.058754e-015, -2.275739e-014, -6.270408e-012, -2.284196e-011,
  5.412204e-014, -2.790928e-014, 4.307576e-011, 5.404352e-011,
  -2.930355e-014, -2.250143e-014, -5.175678e-011, -7.606966e-011,
  2.007857e-014, -1.413994e-014, 7.325576e-012, 1.590554e-012,
  3.35354e-015, -1.620913e-014, -2.361145e-011, -3.154579e-011,
  1.191187e-014, -8.104952e-015, -1.098694e-011, -2.738625e-011,
  1.774405e-014, 1.0126e-014, 3.339456e-011, 3.762361e-011,
  2.199571e-014, 1.249381e-014, 7.28291e-012, 4.413761e-011,
  6.378783e-015, -3.096442e-014, 3.321353e-011, 4.733904e-011,
  6.515428e-015, -4.611836e-016, 5.010985e-011, 5.99363e-011,
  8.820193e-015, -9.809757e-016, -2.893539e-011, -6.326831e-011,
  1.217663e-015, -2.559953e-014, -3.099798e-011, -1.931932e-011,
  1.592191e-014, -1.479299e-014, -5.445614e-011, -8.845926e-011,
  3.854323e-015, -8.647743e-015, -4.66026e-011, -3.206333e-011,
  7.054443e-016, -4.206136e-014, -6.184503e-011, -8.220928e-011,
  1.777139e-014, -4.098557e-015, 3.829837e-011, 3.303122e-011,
  1.020828e-014, -2.301265e-014, -5.943634e-011, -8.380534e-011,
  2.149131e-014, 6.258643e-015, -1.544504e-011, -1.533262e-011,
  4.311981e-015, 2.422642e-015, -2.541594e-011, -1.906312e-011,
  3.047191e-014, -5.577755e-014, 4.101881e-011, 5.461211e-011,
  2.554788e-014, -4.216801e-015, -3.023879e-011, -8.796908e-011,
  3.259659e-014, 3.72429e-014, -5.241071e-011, -6.75017e-011,
  1.969193e-014, -1.686731e-014, 4.685536e-011, 9.938902e-011,
  -3.731062e-015, -3.969444e-014, 3.54284e-013, 1.888503e-011,
  2.768888e-014, -7.785315e-015, -6.559811e-011, -8.245912e-011,
  -1.200366e-015, 4.246955e-014, 2.412792e-011, 2.138223e-012,
  1.454605e-014, 1.573344e-014, 2.287055e-011, 4.492829e-011,
  2.39591e-014, 6.239782e-016, 8.838385e-012, 5.841169e-012,
  2.367881e-014, 1.633148e-016, -2.180267e-012, 1.24838e-011,
  1.968358e-014, 9.096031e-016, -1.65239e-012, -4.0948e-012,
  3.853182e-014, -3.289275e-015, 4.852412e-011, 4.12934e-011,
  2.381247e-014, 2.333657e-015, 2.001504e-012, 4.140696e-012,
  8.824756e-014, -9.445658e-015, -3.043558e-012, 6.643816e-012,
  2.025579e-014, 1.443991e-015, 9.088426e-012, 1.406487e-011,
  2.91678e-014, 1.391196e-015, 1.252007e-011, 2.710273e-011,
  2.378609e-014, 3.936233e-015, -3.642622e-013, -2.551853e-013,
  3.010136e-014, 2.149886e-015, -4.13538e-012, 1.359022e-011,
  2.742543e-014, 3.698581e-015, 4.222846e-013, -1.018311e-011,
  3.11049e-014, 1.676228e-015, -2.113734e-011, 2.547656e-012,
  9.906642e-015, 7.688343e-015, -6.385069e-012, -4.891684e-012,
  1.048185e-013, -7.654843e-015, -5.382085e-012, 1.039035e-011,
  2.997079e-014, -1.151571e-015, -4.44435e-012, -5.370249e-012,
  3.075982e-014, 3.138459e-015, -2.869637e-012, 8.143854e-012,
  4.111596e-014, 5.617374e-016, 1.224134e-011, 5.508127e-012,
  2.394849e-014, 6.221156e-015, 1.062731e-011, 2.216181e-011,
  4.39197e-014, 4.384296e-014, 6.329355e-012, 2.554342e-012,
  5.506629e-015, -1.064803e-013, -3.620324e-012, 1.228901e-011,
  7.09447e-014, -3.753566e-015, 4.14561e-012, 1.860301e-012,
  8.799358e-014, -7.602634e-015, 8.917968e-013, 1.608577e-011,
  3.363574e-014, -5.155053e-016, -1.78335e-012, -4.577512e-012,
  3.938744e-014, -4.755637e-016, 5.341051e-012, 2.054361e-011,
  3.382015e-014, -1.321822e-015, 7.09916e-012, 5.801971e-013,
  3.886495e-014, 5.152496e-015, 5.083385e-012, 1.667998e-011,
  2.920031e-014, 3.298071e-015, 7.97328e-013, -1.861841e-012,
  3.864764e-014, 3.363072e-015, 2.376251e-012, 1.716764e-011,
  3.343222e-014, 1.814588e-015, 3.754227e-012, 3.023517e-012,
  3.713898e-014, 1.647274e-015, 6.303852e-012, 2.045908e-011,
  3.476463e-014, 2.936412e-015, 2.758394e-012, 1.3682e-012,
  3.993289e-014, 1.796653e-015, -5.33939e-012, 1.333842e-011,
  3.4409e-014, 3.263044e-015, -6.826902e-012, -1.222109e-011,
  3.985841e-014, 2.73724e-015, 1.76316e-012, 1.965628e-011,
  3.694826e-014, 1.948621e-015, -2.964546e-013, -1.093623e-012,
  3.822315e-014, 1.697433e-015, 5.01181e-012, 2.239213e-011,
  3.954082e-014, -1.385002e-015, 1.930653e-014, -1.637681e-013,
  3.948431e-014, -4.253512e-016, 4.796839e-012, 2.476314e-011,
  3.696568e-014, 5.202337e-016, 6.846006e-012, 2.528152e-012,
  4.009378e-014, 1.434794e-015, 2.559622e-013, 2.051726e-011,
  4.05448e-014, 8.67767e-016, 2.557563e-012, -2.141389e-012,
  4.591977e-014, 1.546448e-015, -8.255264e-013, 2.353736e-011,
  4.131514e-014, 2.299456e-015, -6.267921e-012, -6.836491e-012,
  4.646921e-014, 3.767989e-017, -5.516968e-012, 1.796994e-011,
  3.813618e-014, 1.278468e-015, -4.908759e-012, -7.238436e-012,
  5.063675e-014, -9.007631e-016, -4.673512e-012, 1.838045e-011,
  -3.962618e-014, 1.191664e-014, -5.693572e-012, -5.260691e-012,
  4.712042e-014, -1.465514e-015, 2.567073e-012, 2.165439e-011,
  4.032994e-014, -2.544718e-015, -3.890513e-012, -3.180641e-012,
  4.587521e-014, -1.692598e-014, 1.05152e-011, 3.218524e-011,
  4.369445e-014, -6.236521e-015, 3.037466e-012, 1.457497e-012,
  5.055546e-014, -9.43294e-015, 4.864054e-012, 2.342425e-011,
  4.421558e-014, -1.963356e-015, 4.434013e-013, -1.313477e-012,
  4.881817e-014, -7.586227e-015, -3.418598e-012, 1.262075e-011,
  9.931169e-015, 2.95612e-015, 5.811858e-012, 1.143654e-011,
  1.215209e-013, -1.86624e-014, -2.12298e-011, 2.021306e-012,
  4.809618e-014, -3.042587e-015, -7.175845e-013, -1.385524e-012,
  5.734365e-014, -3.679144e-015, -6.888042e-013, 1.805551e-011,
  5.238994e-014, -3.075966e-015, -8.095222e-013, 3.218001e-012,
  4.987674e-014, -8.593799e-015, 4.792886e-012, 2.244283e-011,
  5.310838e-014, -7.549849e-015, -4.466914e-012, -5.420821e-012,
  5.773764e-014, -6.67996e-015, -1.486192e-013, 2.525797e-011,
  5.429225e-014, -5.613619e-015, 1.766892e-012, -6.166542e-011,
  6.047444e-014, -5.464631e-015, 8.56786e-012, 6.015117e-011,
  5.420182e-014, -5.500582e-015, 5.635961e-012, -1.381837e-012,
  5.575425e-014, -3.491585e-015, 3.976685e-012, 2.71504e-011,
  7.131235e-014, -6.877713e-015, -2.087766e-012, -1.994213e-012,
  5.577378e-014, -1.959447e-015, 3.846334e-012, 2.906003e-011,
  6.092279e-014, -3.218611e-015, -7.052805e-012, -4.587713e-012,
  6.578411e-014, 1.12222e-015, 5.38056e-013, 2.87309e-011,
  4.970662e-014, -3.498854e-015, 3.453295e-012, 6.04414e-012,
  3.11521e-014, -6.631743e-016, 2.815227e-012, 3.235754e-011,
  4.285063e-014, -5.329205e-015, 3.956707e-012, 1.4615e-012,
  2.498422e-014, -8.437275e-016, 2.834131e-012, 2.981098e-011,
  6.40939e-014, -1.020823e-014, -3.708785e-012, -4.850898e-012,
  7.250021e-014, -6.820041e-015, 5.411289e-012, 3.312281e-011,
  5.879577e-014, -4.871245e-015, -3.809382e-012, -3.584112e-012,
  7.699113e-014, -8.617643e-015, -4.298183e-013, 2.773552e-011,
  6.320283e-014, -2.397778e-015, 1.016865e-012, 4.815324e-013,
  6.352267e-014, -6.453509e-016, -3.336217e-012, 2.870387e-011,
  1.613012e-014, 7.746231e-015, -2.991697e-012, -5.437129e-012,
  -3.075289e-015, 1.474021e-014, 1.113635e-012, 3.356535e-011,
  6.766743e-014, 2.373141e-015, -2.313344e-012, -2.187258e-012,
  7.891733e-014, 2.637478e-015, -4.185625e-012, 3.007103e-011,
  7.443566e-014, 1.584118e-015, 1.018284e-012, -9.871246e-013,
  8.266171e-014, 5.623293e-016, -2.849396e-012, 3.531356e-011,
  7.463212e-014, 2.302659e-015, -2.331894e-013, -8.968411e-014,
  8.069135e-014, 2.473315e-015, -4.177358e-012, 3.534375e-011,
  1.592122e-015, 1.627754e-014, 4.567879e-012, -2.137106e-012,
  6.69111e-014, 9.825324e-015, -3.339315e-012, 3.631213e-011,
  8.262361e-014, 5.385462e-015, -2.228909e-012, -1.938512e-013,
  8.970303e-014, 7.168562e-015, -2.596668e-012, 4.254284e-011,
  8.797931e-014, 1.128103e-014, 8.421224e-013, 4.481718e-012,
  9.499502e-014, 8.656821e-015, -1.425103e-012, 4.86851e-011,
  8.602256e-014, 1.698129e-014, 3.164713e-012, 1.318129e-012,
  9.666287e-014, 1.393507e-014, -3.748542e-013, 4.66303e-011,
  9.423688e-014, 4.473307e-014, 3.495246e-012, 6.539443e-014,
  2.608432e-014, 1.71739e-014, -3.767426e-013, 4.95521e-011,
  9.280556e-014, 1.613051e-014, 1.202767e-011, 4.207723e-012,
  9.515653e-014, 2.269244e-014, 9.63217e-012, 6.139513e-011,
  9.476153e-014, 9.162782e-015, 4.635444e-012, 1.869496e-012,
  1.073453e-013, 2.28912e-014, -1.248422e-011, 4.59618e-011,
  1.013274e-013, 1.430461e-014, 2.441928e-012, -3.217832e-012,
  1.115851e-013, 1.633957e-014, -7.268303e-012, 5.27823e-011,
  1.154418e-013, 8.6986e-015, -2.371007e-012, -4.466411e-012,
  7.318863e-014, 2.109869e-014, -8.97317e-012, 5.209654e-011,
  1.128949e-013, 6.86769e-015, -9.614675e-012, -7.075331e-012,
  9.01766e-014, 1.334253e-014, -7.479378e-012, 5.381946e-011,
  1.146269e-013, 8.889391e-015, -2.99315e-012, -3.916597e-012,
  1.244958e-013, 1.111285e-014, -4.978688e-012, 5.55316e-011,
  1.2006e-013, 4.711987e-015, -2.415207e-012, -6.666036e-012,
  1.34677e-013, 6.01155e-015, -5.363582e-012, 5.523344e-011,
  1.094285e-013, 6.16032e-015, 1.416636e-012, -7.806093e-013,
  1.246631e-013, 4.425554e-015, -1.178143e-011, 5.430062e-011,
  8.502241e-014, 1.164298e-014, 3.935444e-012, 7.202354e-012,
  1.057696e-013, 9.065628e-015, 1.759581e-012, 6.802955e-011,
  1.335674e-013, -1.1232e-015, -3.556728e-012, -3.523715e-012,
  1.541964e-013, -7.182892e-016, 9.137983e-013, 6.782159e-011,
  1.432116e-013, -2.226504e-015, -1.96155e-013, -5.238609e-012,
  1.63455e-013, -4.330715e-016, 4.143787e-012, 7.252443e-011,
  1.464268e-013, -5.280201e-015, 2.46488e-012, -4.39083e-012,
  1.711606e-013, -5.984067e-015, 4.18149e-012, 7.446593e-011,
  1.541753e-013, -7.025692e-015, 2.682753e-012, -1.682049e-012,
  1.765936e-013, -1.071148e-014, 3.536922e-012, 7.614175e-011,
  1.612384e-013, -7.917125e-015, -1.296573e-012, -3.06837e-012,
  1.835481e-013, -1.230357e-014, 5.559722e-012, 7.967834e-011,
  1.655961e-013, -8.844837e-015, 9.056278e-013, -5.514939e-012,
  1.928933e-013, -1.107584e-014, 7.529086e-012, 8.328539e-011,
  1.751578e-013, -1.050644e-014, 8.520173e-012, -8.228327e-013,
  2.081348e-013, -1.059872e-014, 3.740582e-012, 8.499286e-011,
  2.558903e-013, -2.096687e-014, -7.163058e-013, -6.382259e-012,
  1.919049e-013, -1.011959e-014, 4.759694e-012, 8.888551e-011,
  1.913789e-013, -1.035799e-014, -1.464915e-012, -4.388447e-012,
  2.231275e-013, -1.673302e-014, 3.871199e-012, 9.037301e-011,
  2.029816e-013, -1.666866e-014, -8.225426e-012, -1.260636e-011,
  2.407145e-013, -1.201592e-014, 1.016561e-011, 1.049697e-010,
  2.094596e-013, -1.684858e-014, -1.542339e-012, -1.408341e-011,
  2.526702e-013, -1.253033e-014, 1.7888e-011, 1.193886e-010,
  2.826465e-013, -1.975946e-014, -2.610442e-012, -9.737065e-012,
  2.534626e-013, -8.729627e-015, 2.346456e-012, 1.085563e-010,
  2.572855e-013, -1.417569e-014, -1.499627e-012, -9.522959e-012,
  2.727656e-013, -8.772448e-015, 7.496621e-012, 1.156983e-010,
  2.533896e-013, -8.545996e-015, -1.928269e-011, -2.461737e-011,
  2.946712e-013, -1.306354e-014, 2.296255e-011, 1.34693e-010,
  2.626129e-013, -1.239827e-014, -1.882954e-012, -1.136814e-011,
  3.090809e-013, -1.646214e-014, 3.076076e-012, 1.202059e-010,
  2.955465e-013, -1.954874e-014, 5.140917e-013, -1.248166e-011,
  2.935429e-013, -1.111122e-014, 1.123271e-011, 1.324286e-010,
  3.130523e-013, -1.753323e-014, 1.954131e-012, -1.195604e-011,
  2.969798e-013, -5.470702e-015, 9.222031e-012, 1.372005e-010,
  3.146249e-013, -5.607951e-015, 7.231037e-012, -1.220237e-011,
  3.675655e-013, -5.573353e-015, 2.377475e-012, 1.449411e-010,
  3.366555e-013, -1.055582e-015, 4.512993e-012, -1.570065e-011,
  3.804002e-013, -7.165771e-016, -6.354816e-013, 1.532819e-010,
  3.59673e-013, -6.828211e-015, 3.063094e-012, -2.084462e-011,
  3.984787e-013, -2.802132e-015, 1.898674e-012, 1.601127e-010,
  3.872007e-013, -1.418131e-014, 1.68019e-012, -2.460908e-011,
  4.221945e-013, -1.164979e-014, 1.094487e-011, 1.783825e-010,
  4.098361e-013, -2.175688e-014, 3.076828e-014, -2.880251e-011,
  4.542054e-013, -2.147882e-014, 1.103457e-011, 1.861484e-010,
  4.359999e-013, -1.666733e-014, 5.558349e-013, -3.515372e-011,
  4.769059e-013, -1.724552e-014, 9.646465e-012, 1.92608e-010,
  4.637274e-013, -1.557096e-014, 9.608788e-012, -3.817045e-011,
  5.063441e-013, -7.564941e-015, -1.929469e-012, 2.01117e-010,
  5.468486e-013, -1.412702e-014, 5.091962e-012, -4.132609e-011,
  6.051562e-013, -4.103932e-015, 2.570687e-012, 2.270631e-010,
  5.394342e-013, -6.07684e-015, -3.952654e-012, -5.542451e-011,
  5.627204e-013, -2.969849e-015, -7.508588e-013, 2.352735e-010,
  5.831157e-013, -1.630119e-014, -2.635971e-013, -5.107698e-011,
  5.918622e-013, -1.99834e-014, 1.449399e-011, 2.724503e-010,
  6.266013e-013, -1.721387e-014, -5.295175e-012, -6.742085e-011,
  6.20977e-013, -1.92867e-014, 1.515039e-011, 2.987775e-010,
  7.076169e-013, -3.534471e-014, -2.160844e-012, -6.088871e-011,
  7.115567e-013, -3.564921e-014, 1.435876e-011, 3.204219e-010,
  7.341915e-013, -2.853748e-014, -5.266532e-012, -7.06305e-011,
  6.932694e-013, -3.274624e-014, 1.012669e-011, 3.486325e-010,
  7.773829e-013, -3.614126e-014, -1.375008e-011, -7.670185e-011,
  7.119337e-013, -3.995838e-014, 9.260865e-012, 3.76855e-010,
  8.306787e-013, -5.855212e-014, -3.746307e-012, -6.875437e-011,
  7.446677e-013, -6.698481e-014, -3.414417e-012, 3.98956e-010,
  9.268912e-013, -6.548054e-014, 2.230033e-012, -7.212998e-011,
  7.828946e-013, -5.609356e-014, 2.465434e-011, 4.609865e-010,
  9.564624e-013, -5.071646e-014, 7.396776e-012, -6.322522e-011,
  8.141963e-013, -4.429611e-014, 2.747627e-011, 5.262375e-010,
  9.770793e-013, -3.862641e-014, 1.643191e-011, -5.892746e-011,
  8.509204e-013, -2.943863e-014, 1.24955e-011, 5.717329e-010,
  1.0244e-012, -2.686536e-014, -1.483425e-011, -7.446575e-011,
  8.830037e-013, -2.515186e-014, 3.202778e-014, 6.322416e-010,
  1.066679e-012, -3.521885e-014, -1.355454e-012, -4.681321e-011,
  9.348992e-013, -2.436268e-014, 1.760275e-011, 7.176533e-010,
  1.085581e-012, -3.982624e-014, -8.757715e-012, -3.480059e-011,
  9.976236e-013, -3.868911e-014, 3.120198e-011, 8.09251e-010,
  1.097926e-012, -4.040045e-014, -4.224022e-012, 1.19818e-012,
  1.060163e-012, -4.038612e-014, 3.231689e-011, 8.957398e-010,
  1.100173e-012, -2.871823e-014, 7.866961e-012, 4.993269e-011,
  1.147437e-012, -2.45414e-014, 1.493869e-011, 9.873962e-010,
  1.079685e-012, -2.045483e-014, 4.588984e-012, 1.067443e-010,
  1.255993e-012, -1.748561e-014, 1.622148e-011, 1.096572e-009,
  1.038354e-012, -1.606352e-014, 1.887046e-012, 1.809506e-010,
  1.400378e-012, -1.959565e-014, 1.912729e-011, 1.209566e-009,
  9.671142e-013, -3.659616e-015, 1.210182e-012, 2.770971e-010,
  1.59128e-012, 1.142141e-014, 3.703991e-012, 1.326877e-009,
  8.651501e-013, 1.611309e-014, 4.417956e-012, 4.002868e-010,
  1.848146e-012, 4.205075e-014, -8.848128e-012, 1.447392e-009,
  7.349628e-013, 2.111539e-014, 1.251505e-011, 5.618291e-010,
  2.133233e-012, 5.655218e-014, -1.120276e-012, 1.572079e-009,
  5.180626e-013, 1.553277e-014, -4.389349e-012, 7.215932e-010,
  2.673357e-012, 3.000155e-014, 1.500322e-011, 1.700225e-009,
  3.173615e-013, 1.711924e-014, -3.934207e-011, 9.551064e-010,
  3.276697e-012, 2.568049e-014, -4.395655e-011, 1.746542e-009,
  2.659947e-014, 2.238379e-014, 3.181502e-011, 1.26314e-009,
  4.045048e-012, 2.183885e-014, -7.188359e-011, 1.78978e-009,
  -2.320687e-013, 1.742173e-014, 1.321966e-011, 1.561079e-009,
  5.236026e-012, 8.399714e-015, 7.703436e-013, 1.923851e-009,
  -5.208687e-013, -1.248361e-014, 3.139569e-011, 1.947697e-009,
  6.691058e-012, -8.845449e-014, 2.530284e-011, 1.932795e-009,
  -8.040051e-013, -6.305603e-014, 4.655321e-011, 2.359826e-009,
  8.614238e-012, -2.258755e-013, 5.744749e-011, 1.865246e-009,
  -9.874077e-013, -7.512003e-014, 5.140744e-011, 2.860137e-009,
  1.111235e-011, -2.62239e-013, 6.411506e-011, 1.705239e-009,
  -1.004081e-012, -9.489086e-014, 5.872523e-011, 3.410592e-009,
  1.438476e-011, -3.133422e-013, 5.357143e-011, 1.420855e-009,
  -7.072418e-013, -1.8155e-013, 7.554285e-011, 4.001728e-009,
  1.860723e-011, -4.979788e-013, 7.708332e-011, 9.637966e-010,
  7.179498e-014, -3.726402e-013, 1.197883e-010, 4.622791e-009,
  2.414367e-011, -8.60807e-013, 1.117069e-010, 2.489793e-010,
  1.661316e-012, -6.28954e-013, 1.566671e-010, 5.217187e-009,
  3.127056e-011, -1.259639e-012, 1.455822e-010, -7.694511e-010,
  4.426158e-012, -1.044854e-012, 1.978688e-010, 5.732281e-009,
  4.055686e-011, -1.771563e-012, 1.756403e-010, -2.219003e-009,
  9.06024e-012, -1.570212e-012, 2.249354e-010, 6.075203e-009,
  5.257875e-011, -2.232887e-012, 1.859089e-010, -4.212055e-009,
  1.667452e-011, -2.730931e-012, 2.977956e-010, 6.106738e-009,
  6.81557e-011, -3.325428e-012, 2.630411e-010, -6.889736e-009,
  2.864671e-011, -4.379368e-012, 3.948607e-010, 5.605632e-009,
  8.812391e-011, -4.638429e-012, 3.28414e-010, -1.045346e-008,
  4.801899e-011, -5.766697e-012, 3.840848e-010, 4.216338e-009,
  1.126712e-010, -5.303161e-012, 2.843692e-010, -1.521198e-008,
  7.779682e-011, -8.244797e-012, 3.80231e-010, 1.312617e-009,
  1.472412e-010, -6.066325e-012, 2.976255e-010, -2.150849e-008,
  1.243953e-010, -1.287572e-011, 4.566232e-010, -4.0337e-009,
  1.912833e-010, -7.775877e-012, 4.315784e-010, -2.998346e-008,
  1.983534e-010, -1.762114e-011, 4.740964e-010, -1.349499e-008,
  2.501166e-010, -8.663462e-012, 5.213601e-010, -4.137822e-008,
  3.172505e-010, -2.319778e-011, 4.434809e-010, -2.964905e-008,
  3.282724e-010, -8.886451e-012, 6.113153e-010, -5.651447e-008,
  5.185224e-010, -3.003425e-011, 5.031421e-010, -5.793576e-008,
  4.361e-010, -8.228183e-012, 8.124585e-010, -7.732454e-008,
  8.718369e-010, -3.845081e-011, 1.00093e-009, -1.082621e-007,
  5.867339e-010, -5.374442e-012, 1.468804e-009, -1.060447e-007,
  1.524958e-009, -6.382425e-011, 3.528232e-009, -2.044335e-007,
  7.980933e-010, -4.890577e-013, 3.359911e-009, -1.475703e-007,
  2.712111e-009, -1.225239e-010, 1.092593e-008, -4.068509e-007,
  1.090133e-009, 6.808171e-012, 6.99685e-009, -2.096977e-007,
  3.837684e-009, -2.854886e-010, 3.425277e-008, -8.979687e-007,
  1.370681e-009, 1.871515e-011, 1.390948e-008, -3.085065e-007,
  -1.354109e-009, -5.958798e-010, 1.001795e-007, -2.07053e-006,
  1.272526e-009, 3.2948e-011, 2.575991e-008, -4.556673e-007,
  -1.118746e-008, -6.264737e-010, 1.599135e-007, -3.456848e-006,
  1.295757e-009, 4.867204e-011, 3.131021e-008, -5.728421e-007,
  -1.320539e-008, -6.15937e-010, 1.598122e-007, -3.868394e-006,
  1.367457e-009, 2.681324e-011, 2.657433e-008, -5.979168e-007,
  -1.019099e-008, -1.031712e-009, 1.078504e-007, -3.249596e-006,
  1.524644e-009, -2.940952e-011, 1.807229e-008, -5.182015e-007,
  8.331094e-011, -1.107388e-009, 4.398075e-008, -1.835592e-006,
  1.677142e-009, -2.701568e-011, 1.130192e-008, -3.750882e-007,
  3.907571e-009, -4.485051e-010, 1.498681e-008, -7.958243e-007,
  1.335138e-009, -3.565271e-012, 6.810289e-009, -2.658122e-007,
  2.57194e-009, -9.700524e-011, 4.748618e-009, -3.69516e-007,
  1.003431e-009, 3.885226e-012, 3.165517e-009, -1.895386e-007,
  1.439521e-009, -1.771428e-011, 1.095537e-009, -1.899013e-007,
  7.413736e-010, 3.88059e-013, 1.123592e-009, -1.371209e-007,
  8.279731e-010, -2.012164e-011, 3.826661e-010, -1.021958e-007,
  5.49414e-010, -5.159913e-012, 5.853849e-010, -1.001995e-007,
  4.98466e-010, -2.496216e-011, 4.034514e-010, -5.571796e-008,
  4.139824e-010, -1.013927e-011, 5.36518e-010, -7.412551e-008,
  3.097999e-010, -2.813757e-011, 6.40247e-010, -2.964132e-008,
  3.157378e-010, -1.308128e-011, 7.713896e-010, -5.51489e-008,
  1.954972e-010, -2.213047e-011, 7.586684e-010, -1.429718e-008,
  2.425202e-010, -1.143403e-011, 8.573126e-010, -4.098694e-008,
  1.24612e-010, -1.323994e-011, 6.712655e-010, -5.22816e-009,
  1.882233e-010, -8.071948e-012, 7.655496e-010, -3.040386e-008,
  7.99718e-011, -6.665467e-012, 5.064381e-010, 1.601541e-010,
  1.464893e-010, -4.948297e-012, 6.442926e-010, -2.221816e-008,
  5.038947e-011, -5.236111e-012, 4.838112e-010, 3.172358e-009,
  1.140842e-010, -4.64642e-012, 5.962676e-010, -1.623926e-008,
  3.055618e-011, -3.802111e-012, 4.473423e-010, 4.736766e-009,
  8.988189e-011, -3.796466e-012, 6.075008e-010, -1.161499e-008,
  1.826735e-011, -3.07629e-012, 4.059822e-010, 5.391934e-009,
  7.033048e-011, -3.437048e-012, 6.170169e-010, -8.066789e-009,
  1.037647e-011, -2.034935e-012, 2.774603e-010, 5.462126e-009,
  5.504476e-011, -2.492527e-012, 5.385546e-010, -5.350515e-009,
  5.276586e-012, -1.072866e-012, 1.619948e-010, 5.323076e-009,
  4.302415e-011, -1.184557e-012, 3.590712e-010, -3.329765e-009,
  2.22327e-012, -1.724349e-013, 3.223749e-011, 4.958155e-009,
  3.358955e-011, 6.155174e-014, 1.897377e-010, -1.773063e-009,
  3.990451e-013, -1.132368e-013, 1.862091e-011, 4.493226e-009,
  2.619639e-011, -1.343905e-015, 1.65379e-010, -6.361508e-010,
  -5.942641e-013, -2.535832e-013, 2.507649e-011, 3.923779e-009,
  2.043362e-011, -2.094034e-013, 1.717023e-010, 1.874677e-010,
  -1.068124e-012, -1.985583e-013, 3.533406e-012, 3.441759e-009,
  1.594603e-011, -1.608266e-013, 1.172127e-010, 7.491676e-010,
  -1.163641e-012, -1.150413e-013, 1.521121e-012, 2.936594e-009,
  1.250684e-011, 5.345129e-014, 1.47449e-010, 1.265275e-009,
  -1.097739e-012, -1.044391e-013, -5.350101e-011, 2.366334e-009,
  9.834736e-012, 2.785807e-013, 9.992714e-011, 1.472591e-009,
  -8.359654e-013, -1.46598e-014, -3.55117e-011, 2.050711e-009,
  7.776467e-012, 1.716764e-014, 1.098221e-010, 1.667599e-009,
  -6.361282e-013, 2.951975e-014, 1.861909e-011, 1.8011e-009,
  6.102217e-012, -1.070883e-013, 9.638899e-011, 1.722628e-009,
  -3.912858e-013, -8.668395e-015, -1.836934e-011, 1.411604e-009,
  4.888667e-012, 4.851772e-014, 2.216225e-011, 1.640961e-009,
  -1.352015e-013, -2.947476e-014, -2.095925e-011, 1.143877e-009,
  3.914631e-012, 6.965628e-014, 6.069954e-012, 1.60656e-009,
  9.225822e-014, -2.225634e-014, 8.977143e-012, 9.552867e-010,
  3.173332e-012, 8.715672e-015, 1.801448e-011, 1.566213e-009,
  2.935109e-013, 1.221814e-015, -6.95059e-012, 7.282625e-010,
  2.619984e-012, 2.074809e-014, 1.590057e-011, 1.485936e-009,
  4.603423e-013, -1.181057e-014, -2.643313e-011, 5.493144e-010,
  2.18241e-012, -6.076708e-015, 2.127882e-011, 1.398651e-009,
  5.957815e-013, -3.491832e-014, 6.432982e-012, 4.358441e-010,
  1.848437e-012, -1.768671e-014, 6.732785e-012, 1.283592e-009,
  6.905877e-013, -6.897974e-014, 5.05465e-012, 3.073011e-010,
  1.599982e-012, 4.974974e-014, -2.544937e-011, 1.147066e-009,
  7.818824e-013, 1.670436e-014, -1.163256e-011, 2.140592e-010,
  1.394048e-012, 5.281842e-014, -1.18763e-011, 1.123207e-009,
  8.301082e-013, 5.030054e-014, -2.46754e-012, 1.610331e-010,
  1.241271e-012, 4.8515e-014, -1.581416e-011, 1.036323e-009,
  8.66642e-013, 4.792124e-014, 2.880669e-012, 9.918236e-011,
  1.121746e-012, 4.723191e-014, -2.621009e-011, 9.400636e-010,
  8.940051e-013, 1.032762e-014, 5.236295e-012, 4.382891e-011,
  1.017983e-012, 2.608705e-014, -2.095477e-012, 8.505515e-010,
  8.982114e-013, 4.254079e-015, 1.001875e-012, 1.305123e-011,
  9.515454e-013, -1.313741e-014, 2.068052e-011, 7.848185e-010,
  8.81327e-013, -5.295696e-014, -1.071111e-011, -2.6587e-011,
  8.893864e-013, -7.17e-014, 1.360091e-011, 6.729327e-010,
  8.578702e-013, -5.278743e-014, 2.718512e-011, 1.991623e-011,
  8.304759e-013, -1.062149e-013, 7.960375e-011, 6.833489e-010,
  8.226322e-013, -1.368798e-013, -5.851734e-011, -1.266289e-010,
  7.955609e-013, -2.020228e-014, 5.212415e-011, 5.799482e-010,
  8.157165e-013, 6.292216e-014, -1.814749e-011, -1.117485e-010,
  6.966956e-013, 1.080618e-013, 2.13919e-011, 5.667293e-010,
  7.567647e-013, -7.961736e-014, 1.186704e-010, 1.769719e-010,
  6.827382e-013, -2.382665e-013, -1.110359e-010, 2.586882e-010,
  7.450568e-013, 3.432963e-014, 9.07521e-011, 1.827252e-010,
  6.316565e-013, -3.994529e-013, -3.45436e-011, 3.758651e-010,
  7.007136e-013, -1.053762e-014, 2.239743e-011, -3.257777e-012,
  6.561683e-013, -8.385069e-014, 4.064063e-011, 4.50447e-010,
  7.021286e-013, 1.488263e-013, 2.382557e-011, -2.286436e-012,
  5.738963e-013, -9.361237e-014, 8.250343e-011, 5.124009e-010,
  6.331684e-013, -3.455398e-014, -1.655667e-011, -8.893528e-011,
  6.169151e-013, -1.092763e-015, 3.280759e-012, 3.294904e-010,
  5.944778e-013, -4.966162e-014, 7.338001e-012, -4.372205e-011,
  5.890598e-013, -6.470953e-014, 3.558254e-011, 3.136704e-010,
  5.694645e-013, -3.421785e-015, 4.816043e-011, 2.491942e-011,
  5.592947e-013, -1.324515e-013, 5.802526e-011, 3.307352e-010,
  4.950732e-013, -1.292671e-014, -2.140398e-011, -1.148393e-010,
  5.358172e-013, 5.576432e-014, 2.658897e-011, 2.7125e-010,
  4.682046e-013, -3.554211e-014, -2.131365e-012, -4.098275e-011,
  4.987934e-013, -6.564962e-014, 3.804308e-011, 2.514934e-010,
  4.73811e-013, -7.617759e-015, -3.541397e-011, -1.209793e-010,
  5.033447e-013, 7.775867e-015, 4.666598e-011, 2.556506e-010,
  4.360136e-013, -7.829414e-014, -6.380084e-012, -5.812935e-011,
  4.791876e-013, -3.933812e-014, 9.933806e-012, 1.82185e-010,
  4.318253e-013, 7.277622e-014, -5.924426e-011, -1.665226e-010,
  4.884535e-013, 1.096739e-013, 3.59467e-011, 2.630204e-010,
  3.737357e-013, -7.181313e-014, 8.243299e-012, -1.330153e-011,
  4.323951e-013, -7.804047e-014, -2.593166e-011, 1.267091e-010,
  3.607261e-013, -2.825889e-014, 2.346898e-011, 6.261799e-011,
  3.881297e-013, -2.062642e-013, 6.734245e-012, 1.745617e-010,
  3.411738e-013, -1.014209e-013, 1.507945e-011, -6.868483e-012,
  3.940744e-013, -5.781584e-014, -1.131761e-011, 1.22273e-010,
  3.06307e-013, -1.09556e-013, -8.538048e-011, -1.919421e-010,
  4.055733e-013, 1.409468e-013, -8.346709e-011, -9.243623e-012,
  3.762211e-013, -9.367852e-014, -3.430192e-011, -4.834837e-011,
  3.438535e-013, -5.569482e-014, 3.675731e-011, 1.37426e-010,
  2.902878e-013, 1.600786e-014, 4.61501e-012, 2.644408e-011,
  3.21185e-013, -1.986055e-013, 5.734667e-012, 1.3172e-010,
  2.508517e-013, -1.389412e-013, 2.086648e-011, 2.446196e-011,
  3.163459e-013, -8.239631e-014, 5.806522e-011, 1.301852e-010,
  2.870354e-013, 1.14035e-013, -2.541852e-011, -2.992957e-011,
  3.114207e-013, -8.019022e-014, 1.352821e-010, 3.013131e-010,
  3.118504e-013, -8.707117e-014, 3.529836e-011, 8.203029e-011,
  2.621133e-013, -2.116267e-013, 2.818434e-011, 1.032217e-010,
  2.367852e-013, -3.389458e-014, -1.721309e-012, -6.772539e-012,
  2.764775e-013, -1.039427e-013, 2.660697e-011, 1.178184e-010,
  2.114861e-013, -5.499441e-014, -5.62887e-012, -8.861301e-012,
  2.674493e-013, -9.817939e-014, 5.624783e-011, 1.354639e-010,
  2.080378e-013, -3.328041e-014, 1.323873e-011, 1.748642e-011,
  2.469649e-013, -8.19023e-014, 4.554201e-011, 1.242136e-010,
  2.21035e-013, -3.550741e-014, -1.907217e-011, -2.229637e-011,
  1.8423e-013, -5.750656e-014, 2.803445e-011, 1.037047e-010,
  1.879782e-013, -3.863242e-014, -2.226459e-011, -3.386774e-011,
  2.135353e-013, -2.671029e-014, 1.704004e-011, 8.86906e-011,
  1.696165e-013, -4.47787e-014, 1.36738e-013, -5.083131e-012,
  2.153258e-013, -4.521386e-014, 1.261274e-011, 6.975012e-011,
  1.67066e-013, -3.828865e-014, -2.602866e-012, -1.919151e-011,
  2.165853e-013, -2.066035e-014, 1.248105e-011, 7.591183e-011,
  1.518143e-013, -5.023659e-014, 1.203294e-011, 6.767703e-012,
  2.031431e-013, -3.156004e-014, 8.347939e-012, 6.722133e-011,
  1.504799e-013, -3.611788e-014, -1.764256e-011, -2.567835e-011,
  1.902352e-013, -2.882567e-014, 9.357593e-012, 7.181396e-011,
  1.503916e-013, -3.990997e-014, 8.030314e-013, -7.788361e-012,
  1.795814e-013, -1.772883e-014, 1.204524e-011, 7.104781e-011,
  1.430919e-013, -2.565189e-014, 1.421882e-011, 1.691214e-011,
  1.715856e-013, -3.981536e-014, -1.12863e-011, 3.294452e-011,
  1.384401e-013, -3.24614e-015, 1.747149e-011, 2.349104e-011,
  1.810871e-013, -4.585815e-014, 5.721474e-012, 6.591435e-011,
  1.648647e-013, 1.489551e-014, -4.764848e-011, -8.684909e-011,
  2.53291e-013, 5.745436e-014, 4.425009e-012, 8.127543e-011,
  9.65396e-014, -1.926638e-013, -3.464019e-011, -1.011863e-010,
  1.742779e-013, 1.14726e-013, -2.959542e-011, -2.458145e-011,
  1.082197e-013, -8.677648e-014, -2.573215e-011, 2.758704e-011,
  1.201293e-013, -2.096675e-013, 3.066388e-011, 6.809207e-011,
  6.904542e-014, -3.095285e-013, 2.806675e-011, 2.512696e-011,
  1.384129e-013, 9.038737e-015, -5.292125e-011, -1.237951e-010,
  1.676259e-013, 1.400774e-013, 4.399162e-011, 1.286781e-010,
  1.676737e-013, -2.474208e-013, -2.010225e-011, 5.816656e-011,
  1.097953e-013, -8.355049e-014, 7.192212e-011, 1.73538e-010,
  1.142046e-013, -2.227186e-013, 9.9018e-012, -9.248987e-012,
  1.175584e-013, 2.498861e-013, -1.454151e-011, 1.228377e-010,
  6.312156e-014, -5.296224e-013, -5.337012e-011, 6.463383e-011,
  1.223958e-013, 1.408697e-013, -7.782366e-011, -7.057654e-011,
  1.285207e-013, -1.228544e-013, 8.845272e-011, 2.160961e-010,
  1.538171e-013, -8.158331e-014, -2.073244e-011, -6.896137e-013,
  1.307407e-013, -2.280888e-013, -1.747067e-011, 1.416097e-011,
  1.076185e-013, -2.704131e-015, -3.397736e-011, -1.988271e-011,
  1.165244e-013, -1.030387e-013, 5.163281e-011, 1.1435e-010,
  7.220358e-014, 1.692792e-014, -1.791208e-010, -2.698319e-010,
  1.221395e-013, 1.202468e-013, 2.491513e-011, 4.613179e-011,
  9.78929e-014, 6.054827e-014, -6.630545e-011, -8.059588e-011,
  1.1675e-013, -4.131346e-014, 2.721361e-011, 8.769235e-011,
  8.254339e-014, 2.608692e-014, 6.284003e-011, 1.418477e-010,
  1.366182e-013, -2.67045e-013, 7.274564e-011, 1.493107e-010,
  1.183437e-013, 1.673628e-013, -4.591715e-011, -5.483185e-011,
  1.379426e-013, -6.033307e-014, 5.418306e-011, 1.773316e-010,
  3.12583e-014, -2.206281e-013, 4.975101e-011, 1.505777e-011,
  7.409886e-014, -1.267013e-014, -2.158172e-010, -2.720456e-010,
  6.508685e-014, 2.211517e-014, 4.373167e-012, -1.339232e-010,
  1.258519e-013, 3.069012e-013, -1.12163e-010, -8.774051e-011,
  7.123165e-014, -6.537957e-015, -6.664562e-011, -1.204109e-010,
  1.149983e-013, 5.925726e-014, 1.564537e-011, 5.602965e-011,
  9.230102e-014, 6.599764e-014, 7.551715e-011, 1.02831e-010,
  1.303944e-013, -9.614611e-014, 2.562397e-011, 7.218923e-011,
  6.792013e-014, -5.192646e-014, 2.538815e-011, 1.159256e-010,
  4.997146e-014, -1.9594e-013, 1.421061e-012, -3.637329e-012,
  5.725429e-014, -2.366639e-014, 9.130335e-012, 2.133349e-012,
  8.573356e-014, -8.752319e-016, -3.228557e-012, 1.932254e-011,
  7.481322e-014, -4.987964e-014, -2.660016e-011, -3.950034e-011,
  8.940811e-014, -1.880038e-014, -2.222791e-011, -2.133847e-011,
  1.224898e-013, -2.98696e-014, -2.283543e-011, -3.405597e-011,
  1.250334e-013, -3.558732e-014, -2.391136e-011, -1.570408e-011,
  5.509453e-014, -9.364682e-015, -8.696539e-012, -1.943984e-011,
  7.524302e-014, -1.453267e-014, 9.363755e-013, 1.742556e-011,
  6.018382e-014, -1.617569e-014, -5.407863e-012, -9.846469e-012,
  6.736524e-014, -1.638719e-014, 1.497596e-011, 3.247226e-011,
  5.366048e-014, -2.107252e-014, -4.320556e-012, -8.050817e-012,
  7.277202e-014, -2.609601e-014, 1.381386e-011, 3.474851e-011,
  5.265336e-014, -2.166672e-014, 3.972069e-012, 8.982089e-012,
  6.885878e-014, -2.734283e-014, 8.909296e-012, 2.633382e-011,
  5.279908e-014, -2.568417e-014, -4.145874e-012, -1.637582e-012,
  6.361831e-014, -2.333682e-014, 1.370576e-011, 2.756904e-011,
  5.072407e-014, -3.279319e-014, -2.303711e-011, -2.441801e-011,
  5.670403e-014, -2.724466e-014, 9.026692e-012, 1.956954e-011,
  4.958277e-014, -2.434555e-014, -1.511637e-011, -1.519385e-011,
  4.176224e-014, -3.043466e-014, 1.480788e-011, 2.763143e-011,
  2.51802e-014, -1.348212e-014, 3.586675e-013, 5.862035e-012,
  1.00973e-013, -4.937289e-014, 1.56361e-011, 1.996166e-011,
  4.277987e-014, 1.714741e-015, 4.924266e-012, -1.066788e-011,
  8.431363e-014, -1.510042e-014, -6.564083e-012, 6.327607e-012,
  4.85101e-014, 7.050887e-014, -3.730842e-012, 1.00066e-012,
  9.039834e-014, -4.473812e-014, 2.050704e-011, 6.956081e-011,
  3.604807e-014, -1.582986e-014, 3.548277e-012, 1.664418e-011,
  5.886321e-014, -5.079655e-014, -3.16397e-012, 1.336471e-011,
  5.619242e-014, -6.334732e-015, 3.241228e-012, 7.986556e-012,
  7.072094e-014, -3.208097e-014, -1.328338e-011, 3.341357e-012,
  7.680477e-014, -2.108161e-014, 8.92517e-012, 6.889683e-012,
  8.895976e-014, -3.013107e-014, -6.879598e-014, 2.309771e-011,
  2.727494e-014, -3.506079e-014, 1.051214e-011, 1.008876e-011,
  4.947706e-014, -3.730946e-015, -5.332067e-012, -8.294219e-012,
  4.383728e-014, -2.489324e-014, -4.94217e-011, -6.022693e-011,
  5.483337e-014, -1.910614e-014, 5.403122e-011, 7.230871e-011,
  3.288606e-014, -1.912392e-014, -5.792608e-011, -7.437063e-011,
  5.566635e-014, -1.129985e-014, 2.70096e-011, 3.401436e-011,
  4.046419e-014, -1.632859e-014, 1.347131e-010, 1.5924e-010,
  1.562598e-014, 2.316498e-015, 1.084152e-010, 7.330122e-011,
  1.701116e-014, -1.276447e-014, 1.888335e-011, 2.292249e-011,
  2.691946e-014, -5.44442e-015, 4.656617e-011, 3.325272e-011,
  2.772459e-014, -1.420813e-014, -9.910659e-012, -2.47294e-011,
  5.581026e-014, -1.874628e-014, -2.31262e-011, -1.168954e-011,
  6.882156e-014, -4.543151e-015, -7.233736e-011, -5.967311e-011,
  2.118934e-014, -1.843312e-014, 6.034116e-011, 9.957347e-011,
  -6.402165e-015, 1.86446e-014, -6.013912e-011, -7.440697e-011,
  1.230361e-013, -2.279248e-014, 1.011477e-010, 1.503929e-010,
  1.201896e-014, 1.845017e-014, -1.577315e-010, -2.071356e-010,
  7.227432e-014, -6.802154e-015, -2.174693e-011, 1.102258e-011,
  3.313876e-014, -1.889597e-014, -4.345883e-011, -7.540783e-011,
  4.055553e-014, 3.699068e-014, -9.241656e-011, -1.068384e-010,
  4.225042e-014, 9.419848e-015, 7.056253e-012, 1.005453e-011,
  5.792064e-014, -5.584139e-014, 4.466352e-011, 1.01592e-010,
  4.721455e-014, 9.01634e-014, 4.140033e-011, 2.639306e-011,
  1.081079e-013, -4.966964e-014, -7.486126e-011, -1.470968e-011,
  4.972966e-014, 8.196139e-014, -4.522189e-011, -1.868718e-010,
  1.169972e-013, 3.63495e-013, 2.55635e-011, 7.24437e-011,
  3.386513e-014, 5.446729e-014, 7.353311e-011, 4.943902e-011,
  2.451879e-014, -7.34183e-014, -1.496386e-010, -1.481066e-010,
  3.203403e-014, 6.761062e-014, -3.683612e-012, -4.815054e-011,
  4.321235e-014, 1.288109e-013, -1.086901e-010, -1.231292e-010,
  5.40726e-015, -3.995609e-014, -1.462205e-011, -4.303896e-011,
  4.630584e-014, 2.684272e-014, -2.446532e-010, -2.895688e-010,
  3.339017e-014, -2.06857e-015, -2.427791e-010, -2.026166e-010,
  1.785574e-014, 9.540839e-015, 6.819582e-011, 6.379706e-011,
  3.474877e-014, -2.510404e-014, -2.278159e-011, -3.657748e-011,
  4.78104e-014, 1.214176e-013, 8.177894e-011, 9.374936e-011,
  1.939636e-014, 2.081138e-014, -5.689861e-011, -8.191768e-011,
  4.037029e-014, 3.058478e-014, -2.045615e-012, 1.325357e-011,
  9.920766e-015, -7.407769e-015, 2.200309e-012, -3.164071e-012,
  4.601036e-014, -1.86911e-015, 4.401748e-011, 5.292219e-011,
  -3.004233e-014, -1.061083e-014, 4.816963e-011, 5.480661e-011,
  4.940924e-014, -1.977934e-014, 2.492599e-011, 3.728709e-011,
  3.142625e-014, -7.722199e-015, 3.330291e-011, 3.752568e-011,
  2.205028e-014, -1.642838e-014, 2.640224e-011, 3.931754e-011,
  1.789683e-014, -8.221659e-015, 8.065361e-013, 8.479378e-012,
  2.430869e-014, -7.2196e-015, 4.369528e-012, 1.092133e-011,
  1.616534e-014, -1.476996e-014, -6.454679e-011, -6.410212e-011,
  2.849347e-014, -3.12622e-014, -4.213832e-011, -3.930668e-011,
  1.119713e-014, -4.587848e-015, -3.428303e-011, -4.245394e-011,
  1.082512e-013, -4.111108e-014, -8.599576e-012, 2.786414e-012,
  2.758031e-014, -5.519528e-015, -6.805467e-013, -2.783823e-012,
  3.782002e-014, -1.748062e-014, 3.99127e-012, 1.498477e-011,
  1.562305e-014, -3.575196e-014, 4.923584e-011, 5.007509e-011,
  2.511444e-014, -2.352249e-014, -1.111596e-011, -2.621227e-011,
  2.880204e-014, 6.693428e-014, -1.308543e-012, -6.879031e-011,
  5.943738e-014, 1.475889e-013, -3.728872e-011, -9.61907e-012,
  3.018005e-014, 1.92876e-014, -3.948217e-012, 2.173204e-012,
  2.276535e-014, -5.911673e-014, 5.700232e-011, 1.030555e-010,
  3.298026e-014, 1.335468e-014, 9.415239e-011, 1.225267e-010,
  1.406837e-014, -6.96131e-014, 1.826529e-011, 5.03912e-011,
  2.648733e-014, 7.590516e-014, -7.349969e-011, -1.069125e-010,
  2.458354e-014, 5.930451e-014, -1.720266e-011, 2.848333e-011,
  -7.714544e-015, -2.781007e-013, 1.007905e-010, 8.627593e-011,
  1.869129e-014, 4.660171e-014, -8.22434e-012, -9.253728e-011,
  -1.179066e-015, -5.32824e-014, -4.47773e-011, -7.2114e-011,
  4.780165e-014, 5.799131e-014, -6.733186e-012, -2.681347e-011,
  2.874632e-014, 9.299764e-014, -2.354683e-011, -3.671399e-011,
  2.850989e-014, 5.874676e-015, -2.217839e-011, -1.626922e-011,
  2.461444e-014, 3.62922e-014, 1.660162e-011, 1.702166e-011,
  3.150883e-014, -3.083299e-014, -7.531401e-011, -7.581622e-011,
  2.174006e-014, -4.920541e-015, 4.637066e-011, 6.785871e-011,
  2.846756e-015, -1.109063e-014, -2.619031e-011, -3.268038e-011,
  -9.105081e-015, -1.336311e-013, -7.904249e-011, -1.421926e-010,
  3.719355e-014, 1.281901e-013, -2.851787e-013, -5.205414e-011,
  2.453564e-014, 1.221663e-013, -1.885488e-010, -2.059377e-010,
  -1.047873e-014, 5.193054e-014, -2.95747e-011, 7.29822e-011,
  3.22932e-014, -4.231936e-014, -2.358815e-011, 1.065502e-011,
  9.41756e-015, -1.590598e-013, 3.235283e-011, 5.178931e-011,
  2.890828e-014, 3.850379e-014, 5.047988e-011, 6.484933e-011,
  1.291795e-014, -2.11258e-014, 3.089573e-011, 4.843857e-011,
  -1.588296e-015, 5.709395e-014, 5.134372e-011, 4.339491e-011,
  2.423822e-014, 7.192683e-014, 4.604335e-011, 4.948342e-011,
  -5.283671e-014, 1.539498e-015, -1.495563e-011, -2.884206e-011,
  3.407639e-014, -1.037228e-014, 4.112049e-011, 4.985778e-011,
  1.843116e-014, -6.477676e-015, -2.15635e-011, -4.259969e-011,
  2.477522e-014, 2.988206e-014, 5.444578e-011, 5.745579e-011,
  4.335393e-015, -1.107338e-014, 3.277727e-012, 2.736787e-011,
  1.298502e-014, -5.596134e-014, 8.84209e-012, -2.266973e-012,
  1.344048e-014, 1.199261e-014, -7.73761e-011, -6.600639e-011,
  2.24989e-014, -4.89483e-014, 1.08922e-011, 1.659564e-011,
  2.000107e-015, 1.491946e-014, 1.268015e-011, 7.11402e-011,
  -7.683998e-015, -1.888083e-013, 1.12777e-011, 3.607705e-011,
  8.407163e-015, -4.965066e-014, 1.529988e-012, -3.644046e-011,
  3.321748e-014, 1.13246e-013, -4.114645e-011, -5.32602e-011,
  1.975327e-014, -3.182602e-014, 9.994602e-011, 1.169895e-010,
  2.369176e-014, -1.431894e-014, 4.7331e-011, 5.060457e-011,
  -2.117034e-015, -3.375537e-014, 3.328011e-011, 6.481454e-011,
  1.145673e-014, -8.534919e-014, -6.757571e-011, -1.025407e-010,
  -1.6931e-014, -4.397299e-014, 8.018806e-011, 8.219489e-011,
  -4.273587e-014, -4.141007e-014, -8.71261e-011, -1.276212e-010,
  -3.825757e-014, -1.055948e-013, -6.829839e-011, -1.305499e-010,
  -1.823519e-015, 9.449656e-014, 8.039192e-013, -2.984579e-011,
  -2.364409e-014, 1.922887e-014, -1.381426e-010, -2.059057e-010,
  3.747948e-014, 1.47692e-013, -1.432663e-010, -1.181952e-010,
  2.861879e-014, 2.320294e-016, -1.441184e-010, -1.619817e-010,
  2.282464e-014, 1.930584e-014, 1.357513e-010, 1.556961e-010,
  -5.254701e-014, -1.776926e-014, -1.451131e-010, -2.307056e-010,
  2.5396e-014, 1.308367e-013, -3.669077e-011, -4.136781e-011,
  -5.027191e-014, 3.612849e-014, -2.204314e-012, 8.748138e-013,
  9.501903e-015, -4.629496e-014, -5.851638e-011, -4.106993e-011,
  9.038522e-015, 2.794061e-014, -1.375319e-010, -1.478394e-010,
  7.085225e-015, -2.050092e-015, -8.528649e-011, -4.027877e-011,
  3.89882e-014, 1.426114e-013, -8.144926e-011, -1.431714e-010,
  3.195151e-014, 1.387912e-013, -8.319818e-011, -2.133293e-011,
  3.845985e-014, 1.336525e-014, -1.303386e-011, -1.412736e-011,
  3.133027e-014, 1.702223e-014, 2.012401e-010, 2.490096e-010,
  2.11617e-014, -6.280606e-014, 1.056119e-011, 1.740278e-011,
  2.179666e-014, -1.932514e-015, -1.38263e-011, -1.302962e-011,
  3.342255e-014, 7.374553e-015, 1.424961e-011, -4.363467e-012,
  3.4228e-014, -2.0381e-014, 4.650432e-011, 9.785845e-011,
  2.950442e-014, 3.464199e-014, 8.160869e-011, 9.842177e-011,
  9.23032e-015, -6.060315e-014, 8.127007e-011, 1.043175e-010,
  2.290046e-014, -2.49585e-014, 8.57629e-013, -8.746858e-012,
  2.123648e-014, 1.718113e-014, 7.462576e-011, 6.054575e-011,
  1.876745e-014, 1.735339e-014, -2.537393e-011, -4.230414e-011,
  -4.688701e-014, -2.563877e-015, 1.104379e-010, 1.332341e-010,
  1.151691e-014, 2.245927e-014, 2.816761e-011, -3.823292e-012,
  2.887977e-014, 6.546968e-014, 2.296012e-011, 4.600908e-011,
  9.679599e-015, 3.523207e-014, 4.375852e-012, 1.957636e-011,
  1.088718e-014, -1.906509e-014, -4.968827e-011, -2.958726e-011,
  4.470979e-014, 1.216866e-013, 5.024405e-011, 9.276808e-011,
  -5.163335e-016, -6.106934e-014, 4.150638e-012, 5.778674e-011,
  -2.138001e-014, -6.627879e-014, 9.085189e-011, 1.295921e-010,
  -3.167111e-014, -8.388211e-015, 3.059981e-011, 3.721978e-011,
  7.408073e-015, 1.699157e-014, -9.379605e-011, -1.561582e-010,
  2.704224e-014, 2.679287e-014, 2.770345e-011, 7.304492e-011,
  9.643574e-015, -5.37749e-015, -1.654222e-011, -3.379853e-011,
  1.293911e-014, 5.323054e-015, 1.297412e-011, 3.432833e-011,
  -1.043357e-014, 3.057499e-014, -5.601816e-012, 5.019993e-012,
  -5.784598e-015, -4.819266e-014, -1.154207e-011, -1.137068e-011,
  1.114073e-014, -7.056034e-014, 5.023827e-011, 8.970812e-011,
  -7.828118e-015, -5.755005e-014, 6.98898e-011, 6.240724e-011,
  -3.852302e-014, -1.824183e-013, 2.827548e-011, 9.016014e-011,
  -6.4759e-015, -1.373378e-013, -7.274341e-011, -1.352112e-010,
  2.506603e-014, -4.246491e-014, 1.302341e-011, 9.430687e-011,
  -1.204537e-014, -1.463617e-013, -5.904246e-011, -4.134527e-011,
  4.110943e-014, 1.224441e-013, -3.555649e-011, -9.200031e-013,
  -1.226025e-014, -6.619878e-014, -3.23679e-010, -2.786506e-010,
  -1.071361e-015, -6.667692e-014, 1.43895e-010, 1.369959e-010,
  3.467343e-014, 1.117325e-014, 3.235832e-011, 3.193361e-011,
  6.159729e-014, 2.614976e-016, 6.228836e-011, 8.426603e-011,
  2.299959e-014, -5.816373e-014, 8.001858e-011, 1.235758e-010,
  -2.359615e-014, -9.114713e-014, -5.138226e-011, -1.513044e-010,
  8.759828e-014, 3.326334e-013, -2.016113e-010, -2.37611e-010,
  1.257163e-014, -2.482276e-013, 4.800399e-011, 6.849587e-011,
  8.185884e-015, 3.240996e-014, 8.741549e-011, 2.983324e-011,
  -5.468661e-014, -4.875254e-014, 1.704801e-011, -5.662529e-011,
  4.821829e-015, 1.537764e-014, -1.256378e-010, -2.164172e-010,
  1.365082e-014, -1.060345e-015, -4.562696e-012, -6.408458e-012,
  3.782824e-014, 1.607204e-015, 3.82357e-012, 1.295304e-011,
  3.156656e-015, 3.154134e-015, 9.542533e-012, 6.05118e-012,
  3.799462e-014, 1.195797e-015, -3.286358e-011, -8.619827e-012,
  -2.092029e-014, 4.605209e-015, -1.125327e-011, -1.140064e-011,
  7.421583e-014, -3.382663e-015, -5.922415e-012, 3.144734e-012,
  3.373191e-014, 8.406993e-015, -8.20774e-012, -1.664035e-012,
  2.834632e-014, -8.446619e-015, 1.526491e-011, 2.733183e-011,
  2.803238e-014, 4.187533e-015, -2.633156e-013, 1.263732e-012,
  2.739291e-014, 8.56491e-016, 3.325913e-012, 1.635633e-011,
  1.825486e-014, -3.71069e-018, 6.705708e-013, -2.183185e-012,
  2.526618e-014, 1.271203e-015, -1.097011e-011, 1.288058e-011,
  -5.889671e-014, 1.59181e-014, 2.306994e-012, 1.882669e-012,
  4.132241e-014, 2.6707e-015, -1.632118e-012, 1.039246e-011,
  2.650426e-014, 1.255932e-014, 7.238383e-013, 8.992799e-013,
  2.890629e-014, 1.404303e-014, 8.674898e-012, 2.213712e-011,
  -5.631744e-014, 1.418759e-014, -9.132073e-012, -1.468526e-011,
  2.332369e-014, 5.971689e-015, -2.06929e-011, -3.628118e-012,
  -6.996654e-014, -1.054299e-013, -8.248516e-012, -1.423761e-011,
  4.452628e-014, -1.126676e-014, -1.979602e-011, 5.466507e-013,
  -5.333281e-014, 1.452705e-014, 8.602848e-012, 1.657195e-012,
  3.448254e-014, 4.00069e-015, -5.600782e-012, 1.293726e-011,
  2.328296e-014, 4.698458e-015, 2.68881e-012, 8.526723e-013,
  3.367566e-014, 7.003644e-015, -1.910676e-012, 1.369747e-011,
  3.606216e-014, -1.890857e-015, 5.036974e-012, 4.563451e-012,
  3.170023e-014, 2.012225e-015, -6.545642e-012, 6.804972e-012,
  3.566144e-014, -1.881094e-015, -1.238138e-011, -1.518608e-011,
  4.107212e-014, 1.264721e-015, 4.600207e-012, 1.643364e-011,
  2.95071e-014, 3.115004e-015, -4.3669e-012, -5.78414e-012,
  3.415311e-014, 1.215347e-015, 2.293091e-012, 1.336342e-011,
  3.768663e-014, -3.69591e-015, 7.573909e-012, 1.585071e-012,
  2.67014e-014, 3.661004e-015, -2.883997e-012, 5.128913e-012,
  5.013659e-014, -3.348771e-015, 1.311431e-011, 6.629845e-012,
  1.650389e-014, 1.053708e-014, -5.270789e-012, 1.417244e-011,
  3.659868e-014, 2.73828e-015, -3.752467e-012, -2.95638e-012,
  4.608602e-014, 2.79192e-015, 1.896837e-012, 1.747585e-011,
  2.69423e-014, 8.025775e-015, -4.722714e-012, -8.614915e-012,
  4.619445e-014, 2.084946e-015, -2.340007e-013, 1.352416e-011,
  3.214e-014, -2.358094e-015, -1.721272e-012, -3.681251e-012,
  3.259777e-014, 3.7018e-015, -2.832138e-012, 1.071942e-011,
  4.972333e-014, -1.243101e-016, 4.277503e-012, 2.981863e-012,
  2.776945e-014, 2.940527e-015, 1.722748e-011, 2.596936e-011,
  4.570763e-014, 2.692767e-015, 6.638471e-012, 4.841491e-012,
  3.266916e-014, 1.177472e-015, 8.610125e-013, 1.726444e-011,
  4.662744e-014, 1.661422e-015, -1.261859e-011, -9.591976e-012,
  7.555544e-014, -6.661987e-015, -9.244277e-012, 6.194989e-012,
  1.206179e-014, -2.762292e-015, -4.517137e-012, -5.755368e-012,
  1.317124e-013, -9.213384e-015, 2.964233e-012, 1.864216e-011,
  4.526245e-014, -9.987521e-015, 1.932287e-012, -9.288995e-013,
  3.935243e-014, -2.583711e-015, -3.754348e-012, 1.406474e-011,
  3.455852e-014, 6.033116e-016, -5.541034e-012, -5.577789e-012,
  4.740844e-014, -3.64529e-015, 9.164477e-012, 2.240734e-011,
  4.061496e-014, -1.684559e-014, 3.830256e-012, 3.612988e-012,
  4.803777e-014, -4.374673e-015, 7.764468e-012, 2.146111e-011,
  -3.404268e-014, 6.032295e-015, -1.094108e-011, -1.480201e-011,
  1.056255e-013, -1.205046e-014, 9.291038e-013, 1.401461e-011,
  4.157394e-014, 1.05159e-015, -1.051303e-011, -1.051225e-011,
  5.588673e-014, -9.225853e-015, -2.921249e-012, 1.634406e-011,
  4.109372e-014, -3.364542e-015, 1.17891e-011, 6.148476e-012,
  5.125058e-014, -1.036596e-014, 1.137566e-011, 2.437468e-011,
  4.6529e-014, -6.266297e-015, 4.655647e-013, -5.203905e-012,
  5.652654e-014, -9.088875e-015, 8.046964e-012, 2.687859e-011,
  4.739172e-014, -7.349578e-015, 7.501816e-012, -2.51813e-011,
  6.681551e-014, -7.176704e-015, 1.376737e-011, 8.049975e-011,
  5.922107e-014, -3.629608e-015, -1.146096e-012, -3.675038e-012,
  7.580454e-014, -9.987321e-015, 1.799135e-011, 3.993633e-011,
  5.549936e-014, -6.033684e-015, -5.01271e-012, -8.301319e-012,
  6.720622e-014, -5.903046e-015, -2.232073e-012, 1.919369e-011,
  5.735591e-014, -8.200986e-015, 1.004765e-012, -4.342137e-012,
  6.218276e-014, -3.110532e-015, -4.127709e-013, 1.680545e-011,
  1.051983e-013, -1.602449e-014, 4.323652e-013, 2.341672e-012,
  7.538687e-014, -1.972876e-014, 1.039094e-011, 3.221957e-011,
  1.140978e-013, -1.344355e-014, -4.79123e-012, -9.608745e-012,
  6.567389e-014, -9.558331e-015, 6.375141e-012, 2.957402e-011,
  5.693747e-014, -4.056274e-015, -2.929593e-012, -3.015286e-012,
  6.551856e-014, -9.235092e-015, -4.459369e-012, 1.976964e-011,
  4.526163e-014, -1.468965e-015, -3.848234e-012, -2.977773e-012,
  7.051751e-014, -7.591459e-015, 2.073809e-012, 2.501787e-011,
  6.472103e-014, -2.751973e-015, -5.790763e-013, -2.793348e-012,
  8.95323e-014, -4.222192e-015, 3.634248e-012, 3.033943e-011,
  1.136603e-013, -5.928254e-015, -3.543501e-012, -8.236155e-012,
  1.155013e-013, -2.191624e-015, -5.486678e-012, 2.111885e-011,
  7.139532e-014, 1.277893e-015, 7.91383e-012, 3.63435e-012,
  7.20627e-014, 4.863965e-015, -5.450879e-012, 2.636284e-011,
  7.227997e-014, 9.186625e-016, 6.557678e-012, 3.58405e-012,
  7.800829e-014, 4.205972e-015, 2.61836e-012, 3.35273e-011,
  7.287758e-014, 2.50055e-015, -4.789249e-013, -1.861255e-012,
  7.818424e-014, 7.297111e-015, 5.77457e-012, 3.739493e-011,
  8.670654e-014, 2.750007e-015, 6.675406e-013, -2.240743e-012,
  1.678232e-013, -1.17635e-015, -8.219309e-013, 3.516031e-011,
  6.872754e-014, -7.26746e-016, 2.063075e-012, -1.491551e-012,
  9.461761e-014, 3.725613e-015, -4.746497e-012, 2.940213e-011,
  7.214158e-014, 9.086007e-015, -2.533195e-012, -1.017279e-011,
  8.998732e-014, 8.041649e-015, 3.225583e-012, 4.668871e-011,
  7.701999e-014, 1.489768e-014, 3.251801e-012, 9.068312e-013,
  9.076124e-014, 1.808609e-015, -1.18198e-012, 3.862834e-011,
  1.444296e-014, 8.674842e-016, 2.942816e-012, 5.551236e-013,
  1.759455e-014, 3.588409e-015, -1.914668e-011, 2.140052e-011,
  7.445392e-014, 1.449575e-014, 8.406028e-012, -7.439973e-013,
  8.759815e-014, 2.353317e-014, -9.787142e-012, 3.527021e-011,
  9.152842e-014, 1.787823e-014, 3.789025e-013, -3.960708e-012,
  1.022189e-013, 2.28362e-014, -7.568635e-012, 3.782863e-011,
  9.22776e-014, 1.448753e-014, 2.343398e-012, -2.633686e-012,
  1.063764e-013, 1.642152e-014, -6.553521e-012, 4.190564e-011,
  8.783193e-014, 1.475883e-014, -5.587755e-013, -4.990398e-012,
  6.388205e-014, 1.94533e-014, -5.236006e-014, 4.526575e-011,
  8.479161e-014, 1.856918e-014, 3.634245e-012, -6.5842e-012,
  8.142263e-014, 2.092792e-014, -3.158317e-012, 4.698329e-011,
  1.000989e-013, 7.585706e-015, 2.270171e-012, -4.722256e-012,
  1.224009e-013, 9.836753e-015, -4.136729e-012, 4.752791e-011,
  1.065706e-013, 6.003588e-015, -4.902009e-012, -7.576195e-012,
  1.300242e-013, 6.173608e-015, -9.908024e-013, 4.784225e-011,
  1.030847e-013, 8.131572e-015, -1.537933e-012, -6.540947e-012,
  1.077092e-013, 4.732644e-015, -2.742566e-012, 4.710923e-011,
  1.086293e-013, 3.092794e-015, -5.467658e-012, -9.124901e-012,
  7.322268e-014, 8.449854e-015, -8.105315e-012, 4.914679e-011,
  1.215489e-013, -1.931453e-015, -7.083024e-012, -1.083952e-011,
  1.452802e-013, -1.987213e-015, -3.984181e-012, 5.204681e-011,
  1.191927e-013, -2.632007e-015, 2.598398e-014, -4.86576e-012,
  1.501593e-013, -4.091208e-015, 5.91283e-013, 5.547558e-011,
  1.251113e-013, -3.436024e-015, -3.889976e-013, -8.07392e-012,
  1.592135e-013, -6.680302e-015, 3.212266e-012, 6.013628e-011,
  1.317314e-013, -4.614248e-015, 6.350115e-013, -6.851129e-012,
  1.669133e-013, -8.532438e-015, 1.2556e-012, 5.947527e-011,
  1.378715e-013, -6.040762e-015, 1.926288e-012, -4.379426e-012,
  1.692169e-013, -7.96846e-015, 3.886719e-012, 6.623892e-011,
  1.453883e-013, -8.174581e-015, 1.020532e-012, -6.949703e-012,
  1.834952e-013, -1.025082e-014, 5.560215e-012, 7.098617e-011,
  1.492623e-013, -1.018287e-014, -1.10312e-013, -8.570992e-012,
  1.909689e-013, -1.186593e-014, 3.967316e-012, 7.178444e-011,
  7.612581e-014, 1.532145e-014, -4.570459e-012, -1.111382e-011,
  2.296756e-013, -1.212524e-014, 7.072698e-012, 8.175442e-011,
  1.622431e-013, -4.659496e-015, 6.550718e-016, -6.250966e-012,
  2.08978e-013, -1.27539e-014, 5.279422e-012, 7.859818e-011,
  1.633567e-013, -2.578532e-014, 6.093393e-012, -1.441241e-012,
  2.148779e-013, -1.305865e-014, -1.820924e-011, 5.808378e-011,
  1.788261e-013, -3.771693e-014, 2.099002e-011, 8.581476e-012,
  2.291007e-013, -1.869778e-014, -1.010952e-011, 6.148108e-011,
  1.569499e-013, 3.782988e-015, -3.697609e-012, -7.042167e-012,
  1.837347e-013, -3.877273e-015, 7.821609e-013, 8.803454e-011,
  1.808235e-013, -4.337455e-015, -2.425057e-012, -8.166785e-012,
  2.424321e-013, -1.289217e-014, 5.327669e-012, 9.427836e-011,
  2.054e-013, -7.726211e-015, 4.267415e-013, -1.008034e-011,
  2.753124e-013, -1.137256e-014, 2.005902e-012, 9.810237e-011,
  2.253605e-013, -7.508552e-015, 3.656264e-012, -1.016872e-011,
  2.868501e-013, -1.084264e-014, 1.461927e-012, 1.025316e-010,
  2.034979e-013, -2.593382e-015, -3.365237e-012, -1.46064e-011,
  2.903307e-013, -1.171007e-014, 7.17967e-012, 1.101733e-010,
  2.020459e-013, -2.668858e-015, -7.104568e-012, -1.885122e-011,
  3.092587e-013, -6.415004e-015, 3.692518e-012, 1.129002e-010,
  2.699857e-013, -6.673999e-015, -2.451305e-012, -1.446996e-011,
  3.353458e-013, -5.271037e-015, 2.751913e-012, 1.19723e-010,
  2.833011e-013, -2.605498e-015, -8.601821e-013, -1.265087e-011,
  3.605231e-013, -7.288684e-016, 1.409445e-012, 1.252682e-010,
  2.989996e-013, -3.060387e-015, 4.568009e-012, -9.339664e-012,
  3.839039e-013, -7.313044e-015, -1.701455e-012, 1.252167e-010,
  3.194885e-013, -2.219436e-014, -1.306213e-011, -2.032002e-011,
  4.048092e-013, -1.579778e-014, -3.272247e-013, 1.314833e-010,
  3.300037e-013, -2.052937e-014, -2.535153e-012, -2.236266e-011,
  4.223872e-013, -1.79437e-014, 1.736931e-011, 1.550658e-010,
  3.510683e-013, -2.512863e-014, 9.393857e-012, -1.482612e-011,
  4.584825e-013, -1.984399e-014, 2.148168e-011, 1.646461e-010,
  3.614997e-013, -1.968758e-014, -1.885227e-012, -3.463851e-011,
  4.935529e-013, 7.608224e-016, 1.480072e-011, 1.645166e-010,
  4.079172e-013, -1.040859e-014, -6.492539e-012, -4.114841e-011,
  6.165173e-013, -7.444416e-015, 9.629056e-012, 1.808367e-010,
  4.336011e-013, 7.447529e-015, -9.409282e-012, -5.064934e-011,
  5.591512e-013, 2.469344e-015, 6.158651e-012, 1.967209e-010,
  4.672086e-013, 6.339272e-015, 7.908502e-012, -2.987658e-011,
  5.7375e-013, -1.778307e-014, 2.304759e-011, 2.213592e-010,
  5.135307e-013, -1.02773e-014, 1.528593e-011, -3.411807e-011,
  6.15357e-013, -1.10666e-014, 9.085867e-012, 2.213673e-010,
  5.065652e-013, -1.566046e-014, 3.435769e-013, -4.35878e-011,
  6.810799e-013, -2.559538e-014, 1.631578e-011, 2.417747e-010,
  6.157712e-013, -3.011085e-014, 5.946772e-012, -4.531479e-011,
  7.112902e-013, -3.489055e-014, 1.93232e-011, 2.643021e-010,
  6.643625e-013, -3.257289e-014, 4.436457e-012, -5.56105e-011,
  7.330703e-013, -4.145558e-014, 9.790072e-012, 2.793385e-010,
  7.17819e-013, -3.340712e-014, -2.449191e-012, -7.494761e-011,
  7.761489e-013, -4.134978e-014, 1.707126e-011, 3.118445e-010,
  7.260156e-013, -6.44802e-015, -1.343636e-012, -8.395189e-011,
  8.458524e-013, -5.216294e-014, 2.849345e-011, 3.611239e-010,
  8.006702e-013, -4.343496e-014, -8.585697e-012, -9.397634e-011,
  8.82911e-013, -4.188703e-014, 1.48909e-011, 3.780207e-010,
  9.128708e-013, -2.636619e-015, 5.790518e-012, -8.938041e-011,
  9.139991e-013, -1.900023e-014, 2.898965e-011, 4.414637e-010,
  9.618805e-013, -1.061017e-014, -8.318878e-013, -1.041999e-010,
  9.685275e-013, -2.242287e-014, 1.392051e-011, 4.791458e-010,
  1.033132e-012, -1.981325e-014, -1.110337e-011, -1.1855e-010,
  1.019181e-012, -2.696737e-014, 1.068245e-011, 5.30189e-010,
  1.102503e-012, -4.75956e-014, 1.05106e-012, -1.015909e-010,
  1.06207e-012, -3.515032e-014, 2.104062e-011, 6.003228e-010,
  1.158925e-012, -4.121796e-014, -2.709509e-012, -1.0455e-010,
  1.119113e-012, -3.878942e-014, 2.576491e-011, 6.846768e-010,
  1.211826e-012, -2.94322e-014, -6.538048e-012, -1.016991e-010,
  1.190413e-012, -2.740579e-014, 9.529065e-012, 7.591432e-010,
  1.244679e-012, -3.204622e-014, -2.23232e-012, -6.919611e-011,
  1.24597e-012, -2.674156e-014, 1.104353e-011, 8.652639e-010,
  1.264964e-012, -3.05678e-014, -2.418867e-012, -3.716351e-011,
  1.332436e-012, -1.248981e-014, 1.036285e-011, 9.688965e-010,
  1.261053e-012, -9.841965e-015, -9.789286e-013, 1.168184e-011,
  1.44168e-012, 6.801398e-015, 3.509493e-012, 1.097019e-009,
  1.236968e-012, 2.237171e-015, 6.15383e-012, 8.723425e-011,
  1.585023e-012, 4.05379e-014, -3.610571e-012, 1.235688e-009,
  9.421098e-013, 4.620416e-014, 3.628614e-011, 2.149057e-010,
  1.522451e-012, 8.073303e-014, -2.203166e-011, 1.349638e-009,
  9.987071e-013, 8.852743e-015, 3.677025e-011, 3.310215e-010,
  2.021748e-012, 3.380104e-014, 6.382063e-011, 1.5855e-009,
  8.803691e-013, -2.981637e-016, 4.454711e-011, 5.005196e-010,
  2.44408e-012, 8.787714e-015, 1.549841e-011, 1.704028e-009,
  6.961592e-013, 8.974264e-016, 7.376707e-011, 7.768404e-010,
  3.008574e-012, -3.317334e-014, 1.044402e-010, 1.973997e-009,
  3.256981e-013, 6.656509e-015, 3.255226e-012, 9.72038e-010,
  3.64933e-012, 1.636371e-014, 7.031274e-012, 1.983621e-009,
  -4.573575e-014, -1.834443e-014, 2.432748e-011, 1.324032e-009,
  4.635664e-012, -7.028973e-014, 3.58234e-011, 2.105425e-009,
  -4.993178e-013, -3.828675e-014, 1.113003e-011, 1.705004e-009,
  5.977178e-012, -1.666484e-013, 9.460246e-011, 2.209451e-009,
  -9.884988e-013, -4.90543e-014, 3.448371e-011, 2.217397e-009,
  7.783022e-012, -1.858551e-013, 5.730563e-011, 2.173057e-009,
  -1.475097e-012, -5.358557e-014, 5.130715e-011, 2.805655e-009,
  1.027545e-011, -2.393548e-013, 6.763275e-011, 2.10007e-009,
  -1.869177e-012, -8.233727e-014, 6.194871e-011, 3.478519e-009,
  1.360471e-011, -4.067684e-013, 7.565563e-011, 1.862583e-009,
  -2.065664e-012, -1.813347e-013, 9.411975e-011, 4.249085e-009,
  1.814006e-011, -7.460843e-013, 1.214438e-010, 1.41488e-009,
  -1.850687e-012, -3.434575e-013, 1.241723e-010, 5.078153e-009,
  2.418334e-011, -1.128169e-012, 1.525594e-010, 6.799629e-010,
  -9.444711e-013, -6.266775e-013, 1.448209e-010, 5.927067e-009,
  3.232468e-011, -1.639534e-012, 1.602352e-010, -4.859194e-010,
  1.101688e-012, -9.946163e-013, 1.769411e-010, 6.748745e-009,
  4.337182e-011, -2.176629e-012, 1.778074e-010, -2.15891e-009,
  5.482793e-012, -1.87817e-012, 2.792721e-010, 7.461814e-009,
  5.779045e-011, -3.332862e-012, 2.540092e-010, -4.539031e-009,
  1.318027e-011, -3.209878e-012, 3.74968e-010, 7.824059e-009,
  7.703229e-011, -4.82745e-012, 3.162429e-010, -7.855991e-009,
  2.735249e-011, -4.472229e-012, 3.663626e-010, 7.55192e-009,
  1.016626e-010, -5.666132e-012, 2.588891e-010, -1.247991e-008,
  5.048566e-011, -6.896809e-012, 3.633436e-010, 6.092617e-009,
  1.36907e-010, -6.844052e-012, 2.508813e-010, -1.881092e-008,
  8.735258e-011, -1.114224e-011, 4.179825e-010, 2.562755e-009,
  1.830277e-010, -9.113758e-012, 3.380648e-010, -2.759275e-008,
  1.502347e-010, -1.59094e-011, 4.017655e-010, -4.560214e-009,
  2.463667e-010, -1.05825e-011, 4.108738e-010, -3.970922e-008,
  2.553403e-010, -2.177747e-011, 3.521546e-010, -1.779314e-008,
  3.321386e-010, -1.130256e-011, 4.689953e-010, -5.623373e-008,
  4.389508e-010, -2.910337e-011, 3.424664e-010, -4.249803e-008,
  4.531743e-010, -1.103554e-011, 6.784644e-010, -7.945236e-008,
  7.703602e-010, -3.861431e-011, 6.99206e-010, -8.830482e-008,
  6.262308e-010, -8.400141e-012, 1.324632e-009, -1.121926e-007,
  1.397662e-009, -6.591995e-011, 2.898112e-009, -1.790237e-007,
  8.737097e-010, -4.279781e-012, 3.42475e-009, -1.60248e-007,
  2.555823e-009, -1.276693e-010, 9.767955e-009, -3.751447e-007,
  1.219161e-009, 2.980705e-012, 7.577783e-009, -2.332316e-007,
  3.6518e-009, -2.941932e-010, 3.231102e-008, -8.588727e-007,
  1.5541e-009, 1.518587e-011, 1.55913e-008, -3.511856e-007,
  -1.574747e-009, -6.088721e-010, 9.721216e-008, -2.024325e-006,
  1.422687e-009, 3.063326e-011, 2.905768e-008, -5.297407e-007,
  -1.143778e-008, -6.403103e-010, 1.564949e-007, -3.404418e-006,
  1.428101e-009, 5.02961e-011, 3.505467e-008, -6.73128e-007,
  -1.346844e-008, -6.267309e-010, 1.570087e-007, -3.815365e-006,
  1.503946e-009, 2.543572e-011, 2.958449e-008, -7.050095e-007,
  -1.044402e-008, -1.039126e-009, 1.056904e-007, -3.199795e-006,
  1.698295e-009, -4.203197e-011, 1.969276e-008, -6.084704e-007,
  -1.335777e-010, -1.114016e-009, 4.239723e-008, -1.792224e-006,
  1.909075e-009, -3.98026e-011, 1.212306e-008, -4.343602e-007,
  3.728998e-009, -4.529483e-010, 1.392007e-008, -7.589271e-007,
  1.514048e-009, -9.53264e-012, 7.278048e-009, -3.016839e-007,
  2.422623e-009, -9.904454e-011, 4.241815e-009, -3.392366e-007,
  1.118628e-009, 2.315896e-012, 3.273447e-009, -2.104295e-007,
  1.319003e-009, -1.826457e-011, 8.993533e-010, -1.657311e-007,
  8.072329e-010, -2.904796e-013, 1.073609e-009, -1.484348e-007,
  7.319777e-010, -1.965434e-011, 2.954511e-010, -8.307106e-008,
  5.839834e-010, -6.597168e-012, 4.93719e-010, -1.056815e-007,
  4.222867e-010, -2.328742e-011, 3.058379e-010, -4.072793e-008,
  4.289246e-010, -1.209603e-011, 3.935671e-010, -7.597115e-008,
  2.499184e-010, -2.564301e-011, 5.516242e-010, -1.799552e-008,
  3.18725e-010, -1.553971e-011, 6.358442e-010, -5.480294e-008,
  1.488682e-010, -1.975906e-011, 6.466369e-010, -5.384762e-009,
  2.385019e-010, -1.343767e-011, 7.118388e-010, -3.936593e-008,
  8.82985e-011, -1.174614e-011, 5.707584e-010, 1.491126e-009,
  1.79732e-010, -9.460074e-012, 6.58661e-010, -2.810841e-008,
  5.228928e-011, -5.650969e-012, 3.69417e-010, 4.961027e-009,
  1.362324e-010, -5.253462e-012, 5.710476e-010, -1.966341e-008,
  2.942914e-011, -4.116291e-012, 3.821989e-010, 6.692818e-009,
  1.030832e-010, -4.890832e-012, 5.671342e-010, -1.35659e-008,
  1.470326e-011, -2.842803e-012, 3.350829e-010, 7.1589e-009,
  7.89033e-011, -3.903417e-012, 5.711918e-010, -9.059906e-009,
  6.574788e-012, -2.191709e-012, 3.031858e-010, 6.985874e-009,
  6.001766e-011, -3.448045e-012, 5.754986e-010, -5.723889e-009,
  1.897557e-012, -1.486004e-012, 1.889264e-010, 6.404624e-009,
  4.566229e-011, -2.35044e-012, 4.818227e-010, -3.318382e-009,
  -6.907644e-013, -7.397501e-013, 9.287964e-011, 5.79243e-009,
  3.467383e-011, -1.163126e-012, 3.293264e-010, -1.515329e-009,
  -1.860409e-012, -1.830634e-013, -1.215446e-011, 5.056389e-009,
  2.63338e-011, 5.324255e-014, 1.495068e-010, -2.628585e-010,
  -2.242296e-012, -1.247757e-013, -1.051424e-011, 4.332331e-009,
  1.997861e-011, 2.856955e-014, 1.308625e-010, 5.989609e-010,
  -2.173411e-012, -1.771568e-013, 2.416937e-011, 3.652905e-009,
  1.516051e-011, -2.439446e-013, 1.60108e-010, 1.216161e-009,
  -1.879643e-012, -8.986362e-014, 3.507867e-011, 3.041275e-009,
  1.156308e-011, -1.92299e-013, 1.319684e-010, 1.628321e-009,
  -1.472911e-012, 1.447741e-013, -1.841074e-011, 2.443058e-009,
  8.878943e-012, -6.971471e-014, 8.944936e-011, 1.868731e-009,
  -9.731986e-013, 3.288889e-013, -1.026197e-011, 2.005353e-009,
  6.815268e-012, -1.445942e-013, 1.076072e-010, 2.054426e-009,
  -5.329478e-013, -1.12832e-013, -6.384387e-012, 1.523885e-009,
  5.353584e-012, 5.475454e-014, 3.941594e-011, 1.844554e-009,
  -2.516835e-013, -9.326449e-014, -2.115568e-011, 1.173215e-009,
  4.242425e-012, 2.669446e-014, 2.444308e-011, 1.785589e-009,
  1.006247e-013, 3.327974e-014, -1.738402e-011, 9.137224e-010,
  3.396965e-012, 3.835616e-014, 4.724083e-011, 1.765959e-009,
  3.71055e-013, -2.6722e-014, 5.032375e-012, 6.976396e-010,
  2.764216e-012, 3.798209e-014, -4.320361e-012, 1.60993e-009,
  5.829279e-013, -3.38663e-014, -2.795396e-012, 4.983283e-010,
  2.308874e-012, 4.050419e-014, 1.202228e-011, 1.501012e-009,
  7.354413e-013, -3.09541e-014, -1.580776e-011, 3.362904e-010,
  1.962448e-012, 1.924668e-014, 1.819964e-012, 1.375316e-009,
  8.679887e-013, -4.826844e-015, -2.138151e-011, 2.108149e-010,
  1.711323e-012, -1.817278e-015, 6.230222e-012, 1.254581e-009,
  9.456076e-013, -2.55952e-014, -6.510717e-012, 1.353862e-010,
  1.51568e-012, -2.7798e-014, 1.225688e-011, 1.135051e-009,
  9.652826e-013, -1.206559e-013, 1.424625e-011, 8.392913e-011,
  1.373366e-012, -1.398545e-014, -2.891387e-011, 9.594233e-010,
  1.002772e-012, 2.342202e-015, -1.06731e-012, 1.333132e-011,
  1.261681e-012, 3.526221e-014, -2.802059e-011, 8.962053e-010,
  1.01594e-012, 1.669404e-014, -2.383329e-012, -2.609785e-011,
  1.164577e-012, 6.71581e-014, -2.949935e-011, 8.088896e-010,
  1.005048e-012, 4.494067e-014, 1.369217e-011, -4.037283e-011,
  1.085657e-012, 2.316492e-014, -2.63503e-011, 7.398319e-010,
  8.764215e-013, 3.164964e-014, -6.164482e-012, -7.291496e-011,
  1.042171e-012, 1.156069e-014, -2.755942e-011, 6.429954e-010,
  9.300698e-013, -2.917763e-014, -1.039246e-011, -1.088337e-010,
  9.824883e-013, 1.492541e-014, 1.085581e-011, 5.831094e-010,
  8.899027e-013, -9.610512e-014, -2.084278e-011, -9.104391e-011,
  9.202735e-013, -1.492785e-013, 5.130212e-011, 5.34671e-010,
  8.63507e-013, -6.659538e-014, 3.226558e-011, -4.729345e-011,
  8.860756e-013, -8.55626e-014, 5.935845e-011, 5.12447e-010,
  7.549596e-013, -3.428214e-013, -5.208861e-011, -2.93634e-010,
  9.137726e-013, 3.987319e-013, -9.178449e-011, 2.441313e-010,
  7.773836e-013, -4.615562e-014, -3.851888e-012, -1.020833e-010,
  8.940461e-013, 3.884377e-014, 1.023661e-011, 3.715601e-010,
  7.43785e-013, 3.236905e-013, -1.308958e-011, -3.140542e-011,
  7.354885e-013, -3.471521e-013, -2.973585e-011, 3.928121e-010,
  7.12332e-013, 3.111719e-013, -9.979141e-012, -2.695785e-011,
  7.107514e-013, -2.790131e-013, 3.880179e-011, 4.423286e-010,
  6.024278e-013, -2.333631e-014, 9.723826e-012, -3.055774e-011,
  6.846724e-013, -1.042919e-013, -3.066946e-011, 2.442741e-010,
  5.262688e-013, 8.005526e-014, 9.431033e-013, -3.349182e-011,
  6.9514e-013, -1.463086e-013, 4.460056e-011, 3.107447e-010,
  5.171175e-013, -4.329184e-014, 1.238886e-011, -4.461192e-011,
  6.319644e-013, -6.500094e-014, 1.467957e-011, 2.284897e-010,
  4.976335e-013, -3.180158e-014, 9.082969e-012, -3.26268e-011,
  5.989961e-013, -7.397823e-014, 2.587052e-011, 2.295342e-010,
  5.015026e-013, 1.504757e-013, -2.080596e-012, -4.532886e-011,
  5.618413e-013, -7.68468e-014, 4.848863e-011, 2.880944e-010,
  3.673798e-013, -1.727187e-013, -2.743188e-011, -1.19739e-010,
  5.859258e-013, 8.356895e-014, -3.859414e-012, 1.224355e-010,
  3.660893e-013, -5.085675e-014, -9.02818e-012, -5.161815e-011,
  5.358895e-013, -6.15209e-014, 2.95869e-011, 1.780315e-010,
  3.866577e-013, -4.963895e-015, -3.391895e-011, -9.710934e-011,
  4.818958e-013, 4.081811e-014, 2.164954e-011, 1.803968e-010,
  3.64569e-013, -3.456394e-014, -4.094717e-011, -1.013301e-010,
  4.714398e-013, 4.599236e-014, 8.333371e-012, 1.509119e-010,
  3.723529e-013, 1.312927e-013, -7.069541e-011, -1.44022e-010,
  4.667483e-013, 1.283865e-013, 3.794667e-011, 2.195258e-010,
  2.997973e-013, 2.147042e-013, -4.296006e-012, -6.238655e-013,
  4.069761e-013, -1.13077e-013, 3.892111e-011, 2.199386e-010,
  3.432933e-013, 3.528586e-013, 5.456965e-011, 1.026212e-010,
  3.410479e-013, -2.156907e-013, 4.456026e-011, 2.547734e-010,
  2.596155e-013, -1.669679e-013, -5.164806e-011, -1.304204e-010,
  4.183774e-013, 2.002177e-013, -3.054017e-012, 8.202838e-011,
  2.78741e-013, -3.607091e-014, -2.641796e-011, -2.052126e-011,
  3.311639e-013, -1.81915e-013, 1.71919e-010, 3.245353e-010,
  3.622656e-013, -3.107142e-014, 2.70409e-011, 4.957889e-011,
  3.102021e-013, -2.625789e-013, 4.382124e-011, 1.4664e-010,
  2.333725e-013, -7.465765e-014, 2.187986e-011, 6.242409e-011,
  3.030708e-013, -2.644661e-013, 9.370662e-011, 1.905556e-010,
  2.7049e-013, 4.127701e-014, 2.876833e-011, 1.945926e-011,
  2.848205e-013, -8.267021e-014, 9.102298e-011, 2.051393e-010,
  2.445383e-013, 3.691753e-014, 2.873036e-012, 1.845033e-011,
  2.503254e-013, -1.936628e-013, 9.642258e-011, 1.823517e-010,
  2.277397e-013, -4.647983e-016, 9.122271e-013, 7.493835e-012,
  3.176007e-013, -1.467868e-013, 5.120002e-011, 1.291651e-010,
  1.739967e-013, -5.822811e-014, -3.826005e-011, -4.658969e-011,
  2.620404e-013, -8.067425e-014, 2.963548e-011, 9.020362e-011,
  1.842359e-013, -7.78033e-014, 1.861964e-011, 1.998855e-011,
  2.309539e-013, -1.003473e-013, 1.516902e-011, 7.176049e-011,
  1.871572e-013, 6.928368e-014, -3.492555e-012, -3.071359e-012,
  2.300296e-013, -7.066307e-014, 5.684446e-011, 1.564266e-010,
  1.732615e-013, -5.518462e-015, 9.468908e-012, -1.74321e-012,
  2.745867e-013, -5.977509e-014, 1.973247e-011, 9.234362e-011,
  1.477512e-013, -2.921698e-014, -1.179983e-011, -2.130831e-011,
  2.422003e-013, -3.388471e-014, 1.526484e-011, 7.316054e-011,
  1.509252e-013, -1.886351e-014, -1.629299e-011, -2.250708e-011,
  1.971028e-013, -1.271615e-014, 1.738378e-011, 9.249265e-011,
  1.384532e-013, -2.173862e-014, -7.288567e-012, -1.640766e-011,
  1.944265e-013, -2.780633e-014, 1.648342e-011, 7.159592e-011,
  1.467952e-013, -3.529477e-014, -7.023528e-012, -1.176788e-011,
  1.771233e-013, -2.921606e-014, 1.527687e-011, 7.277841e-011,
  1.35011e-013, -1.173524e-014, -2.200474e-011, -4.026932e-011,
  1.725041e-013, 1.212826e-014, 1.271798e-011, 7.114718e-011,
  1.272807e-013, -1.081508e-014, -7.205242e-013, -7.279604e-012,
  1.588736e-013, -8.062509e-015, 1.862783e-011, 6.851077e-011,
  1.294171e-013, 1.571681e-014, 2.541577e-012, -3.011178e-012,
  1.714244e-013, -2.620253e-014, 2.233802e-011, 7.830025e-011,
  1.258777e-013, -2.599907e-014, -1.873615e-011, -4.449201e-011,
  1.683226e-013, 6.283781e-014, 6.615715e-012, 4.895891e-011,
  2.017596e-013, -1.160051e-013, 3.117909e-011, 4.049851e-011,
  1.424755e-013, -1.150352e-013, 3.608957e-011, 6.177836e-011,
  1.166739e-013, 2.291715e-013, 2.403266e-011, 5.493977e-011,
  1.433881e-013, -1.834103e-013, 1.77299e-011, 1.285512e-010,
  8.720172e-014, 1.220421e-014, -1.817138e-010, -3.736169e-010,
  2.546106e-013, 6.338435e-013, -7.058357e-011, 1.296977e-011,
  4.370247e-014, -2.851134e-013, -1.819549e-010, -2.517994e-010,
  1.722788e-013, -1.580018e-013, -1.683485e-011, 1.343628e-011,
  1.572429e-013, -1.210815e-013, 8.135166e-012, -2.673448e-011,
  1.696826e-013, 2.311044e-013, 2.245435e-011, 8.438794e-011,
  1.976549e-013, 7.080811e-013, 1.075836e-010, 2.539087e-010,
  3.51541e-014, -3.718271e-013, 8.052706e-011, 2.964952e-010,
  1.793026e-013, 1.421427e-012, -2.230219e-010, 3.380093e-011,
  -9.51394e-014, -1.446169e-012, 6.095979e-011, 3.474502e-010,
  2.241885e-013, 6.976232e-013, 2.618319e-011, 3.750454e-011,
  6.299625e-014, 5.610881e-014, 9.652017e-011, 2.716964e-010,
  1.389358e-013, -1.20799e-014, 9.524934e-011, 4.327139e-011,
  8.28672e-014, 3.428839e-013, -1.743691e-010, -2.189958e-010,
  6.610841e-014, -3.100674e-013, -1.778943e-011, -4.05328e-011,
  1.392737e-013, 7.938151e-015, -7.719676e-011, -1.314924e-010,
  8.060835e-014, -1.244502e-013, 9.301054e-011, 7.450653e-011,
  1.299967e-013, 8.670207e-015, -2.14084e-010, -2.243837e-010,
  1.154803e-013, -2.062355e-013, 6.25406e-011, 9.960436e-011,
  8.220706e-014, 1.602355e-014, -1.73381e-012, -1.753878e-011,
  -6.731794e-014, -1.760873e-013, -3.115913e-010, -3.392366e-010,
  9.419387e-014, -3.843831e-013, 1.579909e-010, 1.346216e-010,
  7.162112e-014, -3.787346e-014, -1.789646e-010, -5.275858e-011,
  1.352014e-014, -2.427585e-013, 3.187535e-010, 3.370252e-010,
  6.40187e-014, 1.844926e-013, -1.219027e-010, -5.973132e-011,
  -6.062743e-014, -2.437496e-013, 1.641532e-010, 1.512769e-010,
  1.080366e-013, -2.23706e-013, 1.068526e-010, 1.748668e-010,
  5.373044e-014, -3.046311e-013, 2.270347e-010, 2.468543e-010,
  6.094058e-014, -4.523963e-014, 2.638801e-011, -1.879565e-011,
  1.066897e-013, 1.718177e-013, 5.398687e-011, 9.530238e-011,
  2.114227e-014, -5.341191e-014, -5.480509e-012, 3.119733e-012,
  5.512293e-014, -2.371997e-014, 1.651543e-011, 3.27528e-011,
  1.060893e-013, 1.26482e-013, -7.298996e-011, -9.971983e-011,
  8.264238e-014, 9.596515e-014, 5.841387e-011, 1.148986e-010,
  5.572526e-014, 8.833297e-015, -4.625825e-011, -3.835266e-011,
  7.29885e-014, -1.06422e-013, 1.152834e-012, 2.787385e-011,
  4.439176e-014, 5.891561e-015, 1.500726e-011, 1.013537e-011,
  5.427796e-014, -4.185598e-014, -2.069532e-011, 1.801533e-012,
  2.945261e-014, -2.011612e-014, -7.843105e-011, -7.008538e-011,
  1.266318e-014, -5.874497e-014, 1.601235e-011, 4.092737e-011,
  5.836884e-014, -1.555708e-014, -1.162048e-011, -1.99788e-011,
  5.319146e-014, -2.574543e-015, 1.846144e-011, 4.153746e-011,
  4.446205e-014, -8.538882e-015, -8.334552e-012, -1.345835e-011,
  6.310491e-014, -5.404675e-015, 1.174093e-011, 2.457745e-011,
  4.610633e-014, 2.363492e-015, -1.498329e-011, -1.79313e-011,
  4.499658e-014, -1.036831e-014, 1.066339e-011, 2.434342e-011,
  5.298673e-014, -7.51505e-015, 2.098031e-012, 4.855654e-013,
  6.724631e-014, -2.93386e-014, 1.181827e-011, 3.188894e-011,
  6.70726e-014, -3.003542e-014, -1.166745e-011, -1.04619e-011,
  6.829902e-014, -3.703919e-014, 1.289788e-011, 3.13134e-011,
  4.647642e-014, -4.140824e-014, 5.623406e-012, 5.256494e-012,
  5.016149e-014, -3.694982e-014, -2.350884e-012, 6.682818e-012,
  5.39835e-014, -9.362534e-015, -1.3897e-011, -2.135801e-011,
  8.796338e-014, -1.928497e-014, 8.198023e-012, 2.679812e-011,
  7.844647e-014, -4.219015e-014, -4.72412e-012, -1.375585e-011,
  1.0505e-013, -3.706953e-014, 9.596732e-012, 2.600064e-011,
  4.405685e-014, -1.366152e-013, 2.35199e-011, 3.520274e-011,
  5.871691e-014, -5.175663e-014, -3.269346e-011, -4.553586e-011,
  3.685428e-014, 3.366382e-015, 8.51282e-012, 3.064346e-011,
  9.271573e-014, -6.156694e-014, -1.555111e-013, 7.72302e-012,
  1.513871e-014, -2.768521e-014, -3.042561e-011, -2.402704e-011,
  6.85925e-014, -2.992831e-014, -2.137213e-011, -2.577739e-011,
  5.117555e-014, -3.522669e-014, -1.858594e-011, -1.840672e-011,
  8.875339e-014, -2.323382e-014, 1.069816e-011, 1.541131e-011,
  6.138022e-014, 1.19889e-014, -8.658978e-012, -8.833731e-012,
  9.912479e-014, -2.942207e-014, 9.189087e-012, 2.523126e-011,
  2.554313e-016, 5.281774e-014, -1.774729e-011, -1.589325e-011,
  3.506895e-014, -1.65097e-014, -4.761474e-011, -1.667024e-011,
  -2.875685e-014, -2.210759e-014, 3.406464e-011, 5.697254e-012,
  6.630707e-014, 8.5924e-015, -8.167093e-011, -1.067662e-010,
  -2.52506e-014, -1.967355e-014, -3.282493e-011, -6.134484e-011,
  4.533288e-014, 3.208792e-014, -1.267858e-010, -1.436804e-010,
  -9.312465e-014, 3.434151e-014, 2.865913e-011, -2.643649e-011,
  5.201229e-014, -5.110869e-015, -9.72052e-011, -1.314315e-010,
  -3.429659e-014, -5.217778e-015, 8.683988e-012, -2.229236e-011,
  4.898924e-014, -1.484253e-014, -9.523578e-011, -1.078392e-010,
  2.606347e-014, -1.464059e-014, 1.353126e-010, 1.58237e-010,
  3.189889e-014, -1.174587e-014, 2.440493e-011, 2.882758e-011,
  2.830008e-014, -3.806392e-014, -4.455072e-011, 7.922022e-012,
  -7.242258e-014, 8.367697e-015, -2.923952e-010, -3.14445e-010,
  7.509118e-014, -4.142348e-014, -4.627127e-011, 1.138615e-011,
  -1.200714e-013, -1.132248e-015, -3.453253e-010, -3.677741e-010,
  2.579169e-014, 1.411756e-015, -1.912938e-010, -2.28797e-010,
  7.900219e-014, -8.011884e-015, 2.306141e-011, 5.799533e-011,
  5.951067e-014, -5.572804e-014, -9.700808e-011, -1.184526e-010,
  2.064538e-013, 2.662944e-014, 3.294284e-010, 4.368121e-010,
  1.361275e-013, 5.995496e-014, -1.637957e-011, 3.232148e-011,
  3.06392e-014, -9.610493e-014, 1.426821e-010, 2.097909e-010,
  1.149327e-013, 7.680483e-014, 3.813431e-010, 5.441281e-010,
  -5.479398e-014, 1.138756e-013, 6.829912e-010, 7.688288e-010,
  6.986472e-014, -1.362066e-013, 2.365045e-010, 4.290842e-010,
  -5.605465e-014, -3.183658e-013, 1.988171e-010, 2.566834e-010,
  9.103662e-015, 6.988185e-014, 1.216131e-013, -2.783941e-011,
  6.945731e-014, 4.518779e-014, 2.957523e-011, 5.081277e-011,
  1.894947e-014, 7.903883e-014, 6.640071e-011, -9.376395e-011,
  1.6713e-013, 3.374726e-013, 8.086005e-011, 1.259113e-010,
  -1.145489e-013, -2.611519e-013, 5.360574e-011, 4.016539e-011,
  -2.713351e-014, 3.300989e-014, -1.706628e-010, -3.161112e-010,
  -1.133707e-014, -6.888388e-014, -5.335331e-011, -6.171262e-011,
  -3.537786e-014, 1.171328e-013, -3.602377e-011, -8.715877e-011,
  7.767755e-014, 2.709829e-014, 9.565199e-011, 1.182242e-010,
  2.022418e-014, -2.403176e-014, 1.3673e-010, 1.790174e-010,
  8.700728e-015, 1.009493e-013, -4.892421e-012, 2.638706e-012,
  2.868943e-014, -3.473665e-014, 6.813317e-011, 9.919591e-011,
  4.969056e-014, 6.177944e-015, 5.699195e-011, 6.671359e-011,
  5.280909e-014, 3.038377e-015, -1.259968e-011, 5.713771e-012,
  -9.521091e-015, 1.382425e-015, -2.600303e-011, -3.561963e-011,
  9.318449e-014, 1.051849e-014, -5.135065e-012, -9.429524e-013,
  -2.016976e-014, 8.149777e-016, -6.538297e-011, -8.034741e-011,
  5.871379e-014, -2.265852e-014, -2.733717e-011, -3.111881e-011,
  3.242445e-014, -1.5641e-014, 3.490632e-011, 4.151383e-011,
  3.873802e-015, -1.545831e-014, -4.634469e-011, -4.263589e-011,
  -3.459774e-014, -1.61243e-014, 1.90542e-011, 2.960884e-011,
  2.078004e-015, 7.931326e-015, -8.702241e-011, -9.905308e-011,
  -4.310411e-014, -4.706349e-015, 9.391343e-012, 9.942395e-012,
  9.868744e-014, -3.386411e-014, -1.385255e-011, -1.103878e-011,
  1.252448e-014, -3.300251e-014, 1.149867e-011, 2.681008e-012,
  2.742569e-014, -1.941793e-014, -5.085946e-011, -5.01518e-011,
  4.188911e-014, -1.107132e-014, -6.193654e-011, 8.382238e-013,
  -1.87788e-014, -2.141037e-013, 8.043335e-011, 9.379242e-011,
  4.280996e-015, -2.534005e-014, -2.069175e-010, -2.259179e-010,
  5.114603e-014, -1.435722e-013, 9.748264e-011, 1.129545e-010,
  -2.248551e-014, -2.362091e-014, -4.112662e-011, -7.160265e-011,
  5.536053e-014, -4.852841e-014, -2.590416e-011, -4.565412e-011,
  3.168399e-015, -9.247508e-015, 1.262119e-010, 1.574031e-010,
  4.340831e-015, -1.225516e-013, 5.686162e-011, 5.347224e-011,
  -1.921653e-014, -3.780667e-013, 1.303843e-010, 1.466727e-010,
  2.688076e-014, -1.279542e-013, -6.122141e-012, -9.270448e-011,
  -3.705562e-014, -2.62113e-013, 1.097451e-010, 1.383409e-010,
  -2.897953e-014, -3.931252e-014, -7.320328e-011, -1.465951e-010,
  -1.878558e-014, -1.020719e-013, -2.17818e-010, -3.017392e-010,
  6.693586e-014, 7.72715e-014, -1.437165e-010, -1.439566e-010,
  4.937371e-014, -1.670189e-013, -2.110316e-010, -2.265194e-010,
  -3.476747e-015, 1.152335e-013, -1.349789e-010, -1.20292e-010,
  2.673536e-014, 4.501472e-014, -1.047488e-010, -7.746151e-011,
  1.935407e-015, -2.282071e-014, 2.559022e-011, 6.507692e-011,
  -2.006709e-014, 1.05074e-014, -7.288582e-011, -6.827593e-011,
  -1.153493e-014, -2.885443e-014, -7.89723e-011, -8.499222e-011,
  -3.478404e-015, -1.329564e-013, -6.932039e-011, -4.188067e-011,
  1.473584e-015, -8.206214e-014, -2.263387e-013, -2.356084e-011,
  3.551866e-014, 3.304358e-014, 1.312779e-011, 3.759166e-011,
  6.522522e-014, -1.853491e-013, -3.828445e-011, -3.687106e-011,
  -5.70596e-014, -9.97167e-014, 1.185583e-011, -2.138985e-011,
  4.221391e-014, 8.271174e-014, -6.503775e-011, -1.068494e-010,
  -4.55598e-014, -1.297315e-013, 9.008884e-012, -2.413078e-012,
  -2.506274e-014, 8.960409e-014, -1.141966e-010, -1.800175e-010,
  -7.172643e-014, -5.635479e-014, -6.703517e-011, -5.769221e-011,
  4.858696e-014, -1.420618e-013, -2.958078e-011, -5.271683e-011,
  3.808184e-014, -1.705612e-014, -5.538049e-011, -7.51382e-011,
  9.615994e-014, -1.329173e-014, 2.119013e-012, 5.278461e-012,
  9.538917e-016, -8.816523e-014, -5.898738e-011, -4.6238e-011,
  2.255015e-014, -8.166966e-014, 1.733975e-012, -3.904096e-012,
  -9.251343e-015, 7.113146e-015, 7.597226e-011, 1.063441e-010,
  2.784762e-015, -1.625073e-013, -2.48483e-012, 5.996449e-012,
  9.776252e-015, -5.265318e-014, -6.080597e-011, -4.810485e-011,
  6.746732e-014, -8.969934e-014, 2.575558e-011, 1.795445e-011,
  5.698683e-014, 2.024817e-013, 9.775898e-011, 2.286292e-010,
  -5.624044e-014, -5.238361e-013, 1.637771e-010, 2.137805e-010,
  1.214202e-014, 1.439396e-014, 3.538171e-011, 3.873299e-011,
  5.910957e-016, -4.093745e-014, -1.88606e-011, -1.72359e-011,
  1.309466e-014, 4.470682e-015, 1.028114e-011, -1.30642e-011,
  5.084095e-014, 1.60872e-014, 2.539083e-011, 2.885857e-011,
  4.599395e-014, 1.280097e-014, 1.251454e-011, 4.143047e-011,
  -1.794261e-014, -8.513733e-015, 1.464411e-011, 2.713252e-011,
  1.276323e-014, -4.309312e-014, -5.577691e-011, -4.833826e-011,
  -2.573506e-014, -9.558021e-015, -5.159162e-011, -5.180007e-011,
  -4.969879e-014, -1.135606e-013, -3.119194e-011, -7.953023e-011,
  9.803342e-015, 5.553953e-014, -3.65382e-010, -4.097486e-010,
  5.353708e-014, -2.402674e-013, 3.598089e-010, 3.85397e-010,
  6.599095e-014, -1.167663e-014, -2.078452e-010, -2.379106e-010,
  1.20395e-013, -1.505627e-013, 5.959962e-011, 1.365831e-010,
  7.279009e-014, -2.582424e-014, 6.382564e-011, 7.779663e-011,
  4.436861e-014, 2.006188e-014, -5.292856e-011, -3.359818e-011,
  -1.741413e-014, 2.325839e-013, 1.394729e-011, 2.007034e-011,
  -7.684579e-014, 9.984231e-015, -9.622081e-011, -1.264711e-010,
  -5.64832e-014, 1.113963e-014, -8.783992e-011, -1.346324e-010,
  5.11388e-014, -6.247832e-015, -8.108493e-010, -8.543019e-010,
  -1.832442e-013, -1.601587e-014, -5.12119e-010, -6.547922e-010,
  -4.086062e-014, -8.70843e-014, -2.48994e-010, -3.185258e-010,
  3.370515e-014, 6.76122e-014, -1.064544e-010, -1.204451e-010,
  7.169671e-015, 4.822723e-014, -5.741622e-011, -5.41168e-011,
  1.805132e-014, -1.335403e-013, -3.139917e-010, -2.875372e-010,
  5.122913e-015, -6.975972e-015, 1.053754e-010, 5.532436e-011,
  8.077533e-014, -5.426165e-015, -9.45655e-011, -5.428136e-011,
  2.836546e-015, -3.397853e-014, 4.298495e-011, 6.118699e-011,
  -4.803835e-014, 8.166733e-015, -1.029902e-012, -1.628389e-011,
  -2.97568e-014, -4.363484e-014, 4.250812e-011, 4.209172e-011,
  -1.894083e-015, 6.019867e-014, -1.930664e-011, -3.634713e-011,
  8.025828e-014, -2.003487e-014, 2.229011e-014, 1.318232e-010,
  -1.449994e-013, -1.748341e-013, -2.18139e-011, -3.252196e-011,
  3.821215e-014, -1.216644e-014, -4.05423e-011, -4.103666e-012,
  4.227507e-014, -7.63409e-014, 1.126544e-010, 1.388455e-010,
  2.295594e-014, 6.213882e-014, -4.349756e-011, -3.48184e-011,
  5.225957e-015, 2.831977e-014, 4.269193e-011, 6.950698e-011,
  8.262384e-014, 7.130655e-014, 8.861291e-011, 8.058047e-011,
  -5.77635e-014, 1.939053e-013, 3.518003e-011, 7.499497e-011,
  2.86956e-014, -8.38931e-014, -2.320033e-011, -3.126182e-011,
  1.827291e-014, 6.325805e-014, 3.942661e-011, 1.993918e-011,
  -3.878651e-014, 1.422981e-013, 2.189273e-011, 1.944891e-011,
  7.410103e-014, -7.994732e-014, 5.579e-011, 5.655329e-011,
  -4.065882e-014, 2.237046e-014, -1.491468e-011, -3.433301e-011,
  -1.789923e-014, -7.801179e-015, -7.681174e-011, -1.012972e-010,
  -1.766506e-014, 1.593403e-014, -1.591295e-010, -1.823766e-010,
  3.523233e-014, 2.461487e-014, 2.21696e-011, 4.345857e-011,
  -3.860281e-014, -5.45956e-014, -2.52401e-011, -7.968936e-011,
  1.500276e-014, 1.963829e-013, 2.439073e-011, -2.173528e-011,
  1.287943e-013, 1.389727e-013, 1.719332e-010, 1.859331e-010,
  5.439084e-014, 7.223305e-014, 2.079744e-010, 3.009119e-010,
  6.97089e-014, -1.168807e-013, -4.136405e-011, -6.58061e-011,
  6.844841e-014, 2.559073e-013, 1.520632e-010, 1.903221e-010,
  -3.014244e-014, -7.369101e-014, -4.604178e-010, -5.451134e-010,
  5.966685e-014, -2.049786e-014, 2.552598e-011, 2.827825e-011,
  -1.102345e-013, -4.226889e-013, -3.065646e-010, -3.253189e-010,
  -1.229453e-014, -1.603625e-013, -2.757554e-010, -4.130259e-010,
  -8.079745e-014, 9.729504e-014, -3.535555e-010, -4.773237e-010,
  9.136478e-014, 1.347334e-013, 4.220536e-011, 5.343829e-011,
  5.377294e-014, 2.880612e-014, -3.157432e-010, -4.015443e-010,
  1.092942e-013, 1.828058e-013, 3.327744e-010, 4.857576e-010,
  1.807959e-013, 3.168031e-014, 6.360822e-011, 1.551727e-010,
  -4.9839e-014, 2.162721e-014, 1.958066e-010, 2.055804e-010,
  2.503392e-014, 2.06024e-013, 3.323281e-011, 1.356537e-010,
  -2.255172e-013, 4.811652e-014, -3.479231e-010, -5.046442e-010,
  6.059116e-014, -1.408916e-014, 3.689551e-010, 5.620234e-010,
  -6.554094e-014, -2.613843e-013, 4.907694e-011, 5.296988e-011,
  1.965029e-014, 1.215258e-015, -8.364257e-012, -1.00823e-011,
  1.804101e-014, -2.63301e-015, -2.740519e-012, 7.658492e-012,
  -9.28645e-015, 4.933452e-015, -1.194703e-011, -7.978435e-012,
  2.166432e-014, 2.473855e-015, 1.412674e-011, 1.638542e-011,
  -7.697418e-014, 1.752249e-014, 4.425538e-012, 2.954139e-012,
  3.025112e-014, 3.573793e-015, 5.219665e-012, 1.427496e-011,
  8.649076e-015, -5.513965e-015, 3.907993e-012, -3.165158e-012,
  3.079175e-014, 3.100721e-015, 1.24651e-011, 1.583728e-011,
  1.704391e-014, -1.265533e-014, 9.932511e-012, 7.761231e-012,
  2.426158e-014, 2.809646e-015, -2.258629e-012, 1.190917e-013,
  2.082868e-014, -1.723132e-015, 1.876782e-011, 1.662569e-011,
  2.365276e-014, 3.915713e-015, -9.641781e-012, 9.791946e-012,
  -2.974905e-014, 1.066765e-014, 1.310743e-011, 7.434294e-012,
  -4.906918e-014, 8.700559e-015, -8.288565e-012, 2.212352e-012,
  2.007769e-014, 1.410861e-014, -1.366795e-013, -3.501967e-012,
  2.008003e-014, -9.747323e-015, -1.807053e-011, -1.151478e-011,
  -3.728001e-015, 4.678005e-015, 1.278229e-011, 2.528382e-011,
  8.153984e-014, -5.633549e-015, 1.707323e-011, 2.656026e-011,
  2.269221e-015, -6.087244e-014, 1.357857e-011, 2.716003e-011,
  9.69275e-014, 1.118873e-013, 1.652463e-011, 2.780502e-011,
  7.504148e-014, -2.783188e-015, -2.050768e-013, -4.21016e-013,
  -2.486775e-014, 1.66653e-014, -4.122109e-012, 7.302749e-012,
  3.231241e-014, -2.188827e-015, 3.017652e-013, -2.180465e-012,
  1.994765e-014, 8.087789e-015, -7.266618e-012, 3.596516e-012,
  3.063579e-014, 5.102123e-015, -4.265325e-012, -4.159623e-012,
  2.793192e-014, 2.109584e-015, -5.660453e-013, 1.197425e-011,
  1.978091e-014, 3.135502e-015, -8.924609e-012, -9.174741e-012,
  3.671024e-014, 3.564347e-015, 1.38296e-011, 2.78544e-011,
  2.203619e-014, 4.084356e-015, -3.88823e-012, -6.161559e-012,
  4.055471e-014, 3.030277e-015, -3.993771e-013, 1.355446e-011,
  2.784787e-014, 2.752292e-015, 5.1742e-012, 5.510376e-013,
  3.704137e-014, -7.053635e-016, -5.048178e-012, 7.965512e-012,
  2.754054e-014, 5.551523e-015, 2.74864e-011, 3.222311e-011,
  6.503983e-014, -2.785288e-015, -6.783459e-012, 8.444774e-012,
  2.53e-014, 3.486084e-015, 7.372355e-013, -1.699931e-012,
  4.373285e-014, 1.991132e-015, -2.076954e-012, 1.228396e-011,
  2.496995e-014, -3.830655e-015, 2.85325e-012, 3.078264e-012,
  3.756987e-014, 5.924141e-015, -3.395727e-012, 7.944351e-012,
  3.114467e-014, 3.989214e-015, -3.163386e-012, -5.601828e-012,
  2.808773e-014, 1.077303e-015, -1.86121e-012, 1.0427e-011,
  5.098965e-014, -2.132337e-015, 1.274654e-011, 1.106985e-011,
  4.951748e-014, -3.097674e-015, -6.549144e-012, 1.052438e-011,
  4.527757e-014, -6.811603e-015, -3.484161e-012, -2.283067e-012,
  3.666688e-014, -1.193586e-015, -1.627067e-011, -2.40465e-012,
  8.186657e-014, -6.73732e-016, 3.380037e-011, 4.147003e-011,
  6.179247e-014, -3.572545e-015, -1.370311e-011, 4.202341e-012,
  -7.180945e-015, 5.96903e-015, 2.942975e-011, 3.170731e-011,
  1.163901e-013, -4.928584e-015, -5.371122e-012, 5.368732e-012,
  3.609806e-014, -1.091297e-014, 2.101499e-012, -4.02001e-012,
  5.45352e-014, -7.431444e-015, -1.310158e-011, -1.685106e-013,
  3.352825e-014, -1.931346e-015, 2.9012e-012, -1.073515e-012,
  4.725238e-014, -3.404401e-015, 1.869954e-012, 1.540928e-011,
  3.463555e-014, -5.254058e-015, -6.77556e-012, -1.106562e-011,
  4.676862e-014, 6.14447e-015, -2.68949e-012, 1.219321e-011,
  -4.822244e-014, 6.535664e-015, -2.303927e-011, -3.366341e-011,
  7.053449e-014, -5.648468e-015, 2.767527e-011, 4.558227e-011,
  3.511013e-014, -9.959405e-015, -7.409687e-012, -6.888047e-012,
  5.394323e-014, -7.162428e-015, -1.098434e-014, 1.439948e-011,
  4.300976e-014, -4.694705e-015, 7.558012e-012, 5.822522e-012,
  6.399647e-014, -7.938116e-015, 5.436573e-012, 9.530391e-012,
  4.200798e-014, -4.127636e-015, 3.398395e-013, -6.646164e-012,
  5.15066e-014, -4.811253e-015, 5.436185e-014, 1.629686e-011,
  5.32096e-014, -1.073472e-014, -7.679962e-012, -1.205506e-011,
  5.271021e-014, -8.494724e-015, 2.079601e-013, 6.161959e-011,
  3.423155e-014, 4.75781e-017, -1.458086e-012, -5.111354e-012,
  5.660983e-014, -6.136349e-015, 7.321836e-012, 2.496993e-011,
  3.860526e-014, -3.112637e-015, -7.674567e-012, -1.339381e-011,
  8.388428e-014, -8.312075e-015, -4.357178e-012, 1.087965e-011,
  4.912496e-014, 2.451271e-015, -1.174642e-011, -1.315244e-011,
  6.850552e-014, 4.429527e-015, -1.151359e-011, 1.199547e-011,
  1.475351e-014, -4.701393e-015, -2.264238e-012, -1.083184e-012,
  9.972242e-014, -2.465485e-014, 3.516155e-012, 2.224921e-011,
  1.917386e-014, -1.430876e-015, 1.857961e-011, 2.044217e-011,
  1.156151e-013, -2.565715e-014, -1.945241e-011, -5.569745e-012,
  3.555558e-014, -4.101899e-015, -3.501398e-012, -9.066623e-012,
  6.642609e-014, -7.008553e-015, 1.889578e-012, 1.919709e-011,
  5.281512e-014, -4.284388e-015, -3.181527e-012, -8.962252e-012,
  8.067701e-014, -6.968702e-015, 5.056618e-013, 2.063972e-011,
  5.027936e-014, 2.434361e-015, -6.707174e-013, -3.654617e-012,
  5.165337e-014, -1.790951e-015, -3.067091e-012, 2.166312e-011,
  4.313864e-014, 2.411079e-015, -1.140128e-012, -6.704126e-012,
  1.642386e-014, 5.980676e-015, -2.720272e-012, 1.895972e-011,
  6.316533e-014, 2.139038e-015, 3.900053e-012, 1.247897e-013,
  8.047922e-014, -9.779825e-016, 6.691412e-012, 2.743321e-011,
  6.090723e-014, -3.006023e-017, 8.703795e-012, 1.530545e-012,
  7.919573e-014, 4.874012e-015, 6.74218e-012, 3.205435e-011,
  6.009115e-014, 6.58268e-015, -5.317675e-012, -1.282376e-011,
  7.814967e-014, 1.167943e-014, 1.831973e-013, 2.775555e-011,
  1.209745e-013, -4.924441e-015, -1.838731e-012, -7.909387e-012,
  2.580619e-014, 1.827844e-014, -3.770408e-012, 2.865215e-011,
  5.514913e-014, 7.144415e-015, -3.706866e-012, -2.165548e-012,
  7.895715e-014, 1.834523e-016, -4.504844e-012, 2.873292e-011,
  6.364705e-014, 7.347818e-015, 5.062475e-012, 3.923768e-013,
  7.651379e-014, -2.972899e-014, -3.781313e-012, 2.661915e-011,
  6.243922e-014, 9.048987e-015, 3.662043e-012, -2.391404e-012,
  8.433329e-014, 4.346524e-015, -2.457777e-012, 3.276084e-011,
  -3.93532e-014, 3.630716e-014, 1.124732e-012, -7.970978e-012,
  7.0467e-014, 1.136061e-014, 2.228216e-012, 4.39659e-011,
  5.675006e-014, 2.52308e-014, -2.202242e-011, -2.383127e-011,
  9.141687e-014, 2.009748e-014, 5.281146e-012, 4.422855e-011,
  7.847617e-014, 2.041102e-014, -2.43378e-012, -1.421493e-011,
  1.002506e-013, 2.887742e-014, -5.694113e-012, 3.21503e-011,
  7.669713e-014, 1.238903e-014, -8.219757e-013, -8.214305e-012,
  1.018066e-013, 2.119202e-014, -9.141793e-012, 3.073486e-011,
  6.434026e-014, 1.261072e-014, 4.757572e-012, -5.001004e-013,
  7.079779e-014, 2.102736e-014, -6.325508e-012, 3.534351e-011,
  6.297865e-014, 6.92025e-015, 4.870199e-012, -5.269934e-012,
  9.094299e-014, 2.315514e-014, -1.610813e-011, 2.529439e-011,
  8.754419e-014, 5.037106e-015, 4.056324e-012, -3.501311e-012,
  1.182245e-013, 6.094665e-015, 3.03843e-013, 3.853966e-011,
  8.202073e-014, 9.219607e-015, 5.687515e-012, -2.442501e-012,
  1.277135e-013, 7.69637e-015, -1.364391e-013, 4.292371e-011,
  1.072265e-013, 1.437238e-015, 4.800191e-013, -9.465721e-012,
  1.210936e-013, 9.209472e-015, 1.259883e-012, 4.18567e-011,
  1.304e-013, -5.065938e-015, 3.58484e-012, -9.867762e-012,
  8.371136e-014, 2.588016e-014, 1.007523e-014, 4.36884e-011,
  9.672465e-014, 3.7632e-015, -7.885493e-012, -1.739778e-011,
  1.322267e-013, 1.536007e-014, -6.484846e-013, 4.556267e-011,
  1.057697e-013, -1.164678e-015, -1.967275e-013, -5.519975e-012,
  1.395174e-013, -2.358199e-015, -4.106871e-012, 4.542517e-011,
  1.115724e-013, -3.155765e-015, 1.998165e-012, -4.798114e-012,
  1.492434e-013, -5.932398e-015, -7.947311e-014, 5.034501e-011,
  1.17264e-013, -3.163087e-015, 3.048229e-013, -6.377251e-012,
  1.551205e-013, -5.705669e-015, 4.091401e-012, 5.528553e-011,
  1.218004e-013, -5.828043e-015, -2.328976e-013, -7.473329e-012,
  1.615873e-013, -5.588694e-015, 3.07391e-012, 5.600305e-011,
  1.254085e-013, -6.389529e-015, -6.208924e-013, -9.108251e-012,
  1.691874e-013, -7.186024e-015, 2.870518e-012, 5.747401e-011,
  1.312846e-013, -5.227057e-015, -1.118866e-012, -8.025803e-012,
  1.765398e-013, -9.454451e-015, 5.001619e-012, 6.237866e-011,
  2.321456e-013, -3.732504e-014, -9.965227e-013, -9.904265e-012,
  1.488174e-013, -5.338635e-016, -4.280229e-012, 5.512943e-011,
  1.490906e-013, -1.401705e-014, -4.178512e-012, -1.132482e-011,
  1.923743e-013, -8.801713e-015, 2.072111e-012, 6.499244e-011,
  1.514473e-013, -1.597016e-014, -1.29321e-011, -2.558148e-011,
  2.112462e-013, 7.917762e-015, 2.07325e-011, 9.207513e-011,
  1.602626e-013, 1.362612e-015, -8.77528e-012, -2.426185e-011,
  2.236591e-013, 1.22216e-014, 2.785373e-011, 9.866798e-011,
  1.624146e-013, 2.211644e-015, -1.48569e-011, -3.255713e-011,
  3.104248e-013, -1.268639e-014, 1.334353e-011, 8.439652e-011,
  1.798384e-013, -5.684005e-015, -2.138737e-012, -1.310822e-011,
  2.582678e-013, -1.150231e-014, 4.63956e-012, 8.170451e-011,
  1.873168e-013, -8.160159e-015, -1.954322e-011, -2.395968e-011,
  2.454819e-013, -9.0441e-015, -1.547036e-011, 6.751802e-011,
  1.894516e-013, -4.386647e-015, -2.610242e-012, -1.421886e-011,
  2.606888e-013, -1.035999e-014, 6.538499e-012, 8.802996e-011,
  1.86645e-013, -7.452644e-015, 3.741318e-013, -9.867731e-012,
  3.122174e-013, -2.13675e-014, 4.282662e-012, 9.150153e-011,
  1.986028e-013, -6.492596e-015, 4.384819e-012, -9.507612e-012,
  3.487934e-013, -1.72738e-014, 2.162049e-012, 9.69415e-011,
  2.273151e-013, -1.392731e-015, 9.284012e-013, -1.463948e-011,
  3.084815e-013, -7.86266e-015, 2.130385e-012, 1.050317e-010,
  2.425937e-013, 2.818292e-015, 3.723074e-012, -9.460828e-012,
  3.318678e-013, -3.965326e-016, -1.085726e-012, 1.081299e-010,
  2.49778e-013, -1.958467e-015, 2.866403e-012, -9.183427e-012,
  3.641659e-013, -8.432133e-015, 1.166582e-011, 1.267991e-010,
  2.512259e-013, -1.249336e-014, 9.177347e-012, -1.746906e-012,
  3.828045e-013, -3.176908e-014, 2.171717e-011, 1.359537e-010,
  2.708039e-013, -2.052665e-014, -1.012092e-012, -1.797919e-011,
  4.011685e-013, -4.235169e-015, -8.079198e-012, 1.074949e-010,
  2.84163e-013, -2.934555e-014, 5.814357e-012, -2.002197e-011,
  4.412275e-013, 1.169108e-014, -3.458784e-012, 1.147341e-010,
  3.058366e-013, -1.132756e-014, 3.541807e-012, -2.92046e-011,
  4.351038e-013, 1.265023e-014, 5.211464e-012, 1.375688e-010,
  2.767753e-013, -3.428035e-015, 3.795138e-012, -1.825565e-011,
  5.676876e-013, -2.280081e-014, -4.201671e-012, 1.406923e-010,
  3.748903e-013, -2.458801e-015, 1.113093e-011, -9.889158e-012,
  5.3582e-013, -2.170194e-014, 3.650064e-012, 1.645293e-010,
  3.949348e-013, 9.349548e-015, -3.560266e-013, -2.778684e-011,
  5.552683e-013, -1.648683e-014, 1.436977e-011, 1.79925e-010,
  4.156191e-013, -1.213638e-014, -7.217706e-012, -4.19904e-011,
  5.83754e-013, -2.573067e-014, 7.286807e-012, 1.805798e-010,
  4.412183e-013, -1.160869e-014, -1.140206e-011, -4.724357e-011,
  5.652302e-013, -4.305464e-016, 8.239091e-012, 1.964443e-010,
  5.009536e-013, 7.894696e-015, 2.408946e-012, -3.740798e-011,
  6.812656e-013, -4.198138e-014, 8.15164e-012, 2.145679e-010,
  5.575291e-013, 2.845479e-015, -6.15252e-012, -5.390948e-011,
  7.283859e-013, -4.143238e-014, 1.461634e-011, 2.37833e-010,
  6.081215e-013, 6.106767e-015, -8.993748e-012, -6.469815e-011,
  7.753588e-013, -4.961085e-014, 3.874536e-011, 2.825268e-010,
  6.932639e-013, -5.811771e-014, -1.007148e-011, -7.022143e-011,
  7.956083e-013, -5.261143e-014, 2.170209e-011, 2.726634e-010,
  7.448996e-013, -2.604538e-014, 2.088456e-012, -8.00613e-011,
  8.568231e-013, -3.417624e-014, 1.192314e-011, 2.910974e-010,
  7.839316e-013, 1.000224e-014, 1.400938e-011, -7.296714e-011,
  9.326749e-013, -4.163524e-014, 4.397669e-011, 3.719915e-010,
  8.50952e-013, -9.00322e-015, -2.207976e-012, -9.85056e-011,
  9.913966e-013, -3.303466e-014, -3.275527e-012, 3.535592e-010,
  9.270336e-013, -3.373245e-014, -1.000326e-011, -1.244331e-010,
  1.053008e-012, -2.511847e-014, 2.1738e-011, 4.14236e-010,
  1.000283e-012, -6.410955e-014, -1.18385e-011, -1.391361e-010,
  1.117194e-012, -2.339799e-014, 9.508177e-012, 4.384999e-010,
  1.088682e-012, -3.714605e-014, 1.312582e-012, -1.331452e-010,
  1.174188e-012, -4.410596e-014, 6.07829e-012, 5.041852e-010,
  1.175787e-012, -1.882822e-014, 1.041058e-011, -1.269699e-010,
  1.245133e-012, -4.593781e-014, 6.748917e-012, 5.805267e-010,
  1.249066e-012, 1.053176e-015, 3.324957e-012, -1.325998e-010,
  1.305611e-012, -3.342077e-014, 1.970217e-011, 6.821459e-010,
  1.308131e-012, -2.103028e-014, -1.345498e-012, -1.398524e-010,
  1.383888e-012, -1.279764e-014, 1.205895e-011, 7.660182e-010,
  1.363518e-012, -8.214562e-015, 6.722024e-013, -1.224168e-010,
  1.468376e-012, 7.050928e-015, 2.243048e-012, 8.768375e-010,
  1.402631e-012, 1.106781e-014, 4.781067e-012, -8.765716e-011,
  1.567289e-012, 4.847682e-014, -6.12108e-012, 1.006905e-009,
  1.333072e-012, 4.088464e-014, 4.056571e-011, 7.266125e-012,
  1.56448e-012, 5.63564e-014, -2.623178e-011, 1.130021e-009,
  1.370421e-012, 2.289998e-014, 3.599164e-011, 8.499297e-011,
  1.840801e-012, 6.869926e-015, -5.895646e-011, 1.262573e-009,
  1.295269e-012, -1.536908e-014, 1.228722e-011, 1.782398e-010,
  2.082986e-012, 1.163691e-014, 1.880027e-012, 1.469841e-009,
  1.208643e-012, -5.700382e-014, 1.325334e-011, 3.226086e-010,
  2.374411e-012, 3.205295e-014, -1.299306e-010, 1.484983e-009,
  8.983984e-013, 4.43172e-015, 8.970656e-012, 5.172741e-010,
  2.855401e-012, 1.300934e-014, 1.021713e-011, 1.870258e-009,
  5.629215e-013, -4.498916e-014, 2.747035e-011, 8.067575e-010,
  3.502416e-012, -4.683258e-014, 3.613333e-011, 2.070055e-009,
  1.115435e-013, -2.695967e-014, 1.176474e-011, 1.128443e-009,
  4.412636e-012, -1.364542e-013, 7.469784e-011, 2.23992e-009,
  -4.330614e-013, -3.205199e-014, 1.899911e-011, 1.575541e-009,
  5.700163e-012, -1.50692e-013, 6.297996e-011, 2.375102e-009,
  -1.092094e-012, -2.586451e-014, 2.703847e-011, 2.133966e-009,
  7.541768e-012, -2.024511e-013, 5.917253e-011, 2.449586e-009,
  -1.790917e-012, -2.789099e-014, 5.073158e-011, 2.819775e-009,
  1.007682e-011, -3.319023e-013, 7.90886e-011, 2.416819e-009,
  -2.533525e-012, -8.000115e-014, 7.103678e-011, 3.630383e-009,
  1.367108e-011, -6.113253e-013, 1.233369e-010, 2.216298e-009,
  -3.142748e-012, -1.577772e-013, 1.02108e-010, 4.571427e-009,
  1.86373e-011, -9.518797e-013, 1.519283e-010, 1.762493e-009,
  -3.437777e-012, -3.224979e-013, 1.183137e-010, 5.604422e-009,
  2.558391e-011, -1.453257e-012, 1.941294e-010, 9.579133e-010,
  -3.077781e-012, -5.928707e-013, 1.999837e-010, 6.799391e-009,
  3.507651e-011, -1.970434e-012, 1.896894e-010, -3.689861e-010,
  -1.269873e-012, -1.201667e-012, 2.56206e-010, 7.95853e-009,
  4.823176e-011, -3.14879e-012, 2.549442e-010, -2.371912e-009,
  3.065007e-012, -2.189378e-012, 3.563244e-010, 8.988949e-009,
  6.610166e-011, -4.694937e-012, 3.174483e-010, -5.301187e-009,
  1.273699e-011, -3.280127e-012, 3.611639e-010, 9.649476e-009,
  8.983373e-011, -5.712486e-012, 2.616204e-010, -9.564247e-009,
  2.902865e-011, -5.407468e-012, 3.674014e-010, 9.444822e-009,
  1.240455e-010, -7.177032e-012, 2.274313e-010, -1.567027e-008,
  5.883861e-011, -9.391113e-012, 4.208544e-010, 7.598059e-009,
  1.712856e-010, -1.00006e-011, 2.859444e-010, -2.440965e-008,
  1.108967e-010, -1.398631e-011, 3.929413e-010, 2.677766e-009,
  2.367663e-010, -1.196511e-011, 3.208535e-010, -3.680955e-008,
  2.02431e-010, -1.999181e-011, 3.049146e-010, -7.769611e-009,
  3.276704e-010, -1.325216e-011, 3.428504e-010, -5.418434e-008,
  3.685188e-010, -2.776499e-011, 2.607374e-010, -2.879881e-008,
  4.593772e-010, -1.364675e-011, 5.427102e-010, -7.920141e-008,
  6.768986e-010, -3.818135e-011, 4.955787e-010, -6.999833e-008,
  6.505201e-010, -1.142086e-011, 1.196508e-009, -1.151425e-007,
  1.276462e-009, -6.675123e-011, 2.34024e-009, -1.549423e-007,
  9.296555e-010, -8.185628e-012, 3.427023e-009, -1.689211e-007,
  2.401365e-009, -1.311068e-010, 8.648855e-009, -3.440696e-007,
  1.326654e-009, -1.726858e-012, 7.999286e-009, -2.521778e-007,
  3.463341e-009, -3.024301e-010, 3.050519e-008, -8.195245e-007,
  1.71157e-009, 1.003372e-011, 1.70795e-008, -3.883407e-007,
  -1.792888e-009, -6.212793e-010, 9.462871e-008, -1.975036e-006,
  1.538041e-009, 2.610712e-011, 3.211357e-008, -5.975328e-007,
  -1.169296e-008, -6.540969e-010, 1.539494e-007, -3.349875e-006,
  1.511723e-009, 4.879959e-011, 3.874533e-008, -7.671535e-007,
  -1.373047e-008, -6.372041e-010, 1.55171e-007, -3.759028e-006,
  1.593872e-009, 2.203535e-011, 3.258157e-008, -8.04496e-007,
  -1.069618e-008, -1.046239e-009, 1.043668e-007, -3.147345e-006,
  1.830086e-009, -5.720959e-011, 2.136299e-008, -6.914775e-007,
  -3.591119e-010, -1.120085e-009, 4.12642e-008, -1.748201e-006,
  2.110452e-009, -5.493027e-011, 1.288463e-008, -4.871084e-007,
  3.549744e-009, -4.564772e-010, 1.302916e-008, -7.221061e-007,
  1.667301e-009, -1.597341e-011, 7.639675e-009, -3.318164e-007,
  2.277524e-009, -1.009342e-010, 3.81068e-009, -3.099849e-007,
  1.210615e-009, 5.388659e-013, 3.370626e-009, -2.262866e-007,
  1.204417e-009, -1.879231e-011, 7.451487e-010, -1.428651e-007,
  8.548585e-010, -9.863846e-013, 1.05156e-009, -1.558321e-007,
  6.438973e-010, -1.893629e-011, 2.591676e-010, -6.560827e-008,
  6.031149e-010, -7.775694e-012, 4.121221e-010, -1.080383e-007,
  3.549052e-010, -2.129796e-011, 3.258142e-010, -2.749314e-008,
  4.323646e-010, -1.369538e-011, 3.056664e-010, -7.542235e-008,
  1.991693e-010, -2.310249e-011, 5.189403e-010, -8.137825e-009,
  3.132775e-010, -1.754894e-011, 4.892842e-010, -5.274667e-008,
  1.108404e-010, -1.738551e-011, 5.986915e-010, 1.760956e-009,
  2.284487e-010, -1.521602e-011, 5.977417e-010, -3.653985e-008,
  6.044031e-011, -9.880775e-012, 4.814248e-010, 6.518917e-009,
  1.678676e-010, -1.002907e-011, 6.016652e-010, -2.49681e-008,
  3.14515e-011, -4.630564e-012, 3.439316e-010, 8.533653e-009,
  1.237093e-010, -5.589469e-012, 5.05196e-010, -1.666023e-008,
  1.468523e-011, -3.108929e-012, 3.404891e-010, 9.016729e-009,
  9.134527e-011, -4.87334e-012, 5.293964e-010, -1.070968e-008,
  4.229482e-012, -2.004352e-012, 2.870457e-010, 8.582424e-009,
  6.801579e-011, -3.832097e-012, 5.481695e-010, -6.48373e-009,
  -6.259307e-013, -1.510975e-012, 2.310887e-010, 7.727739e-009,
  5.038893e-011, -3.256011e-012, 5.395856e-010, -3.517558e-009,
  -2.858538e-012, -9.433389e-013, 1.543671e-010, 6.711055e-009,
  3.734831e-011, -2.221956e-012, 4.619443e-010, -1.436412e-009,
  -3.675495e-012, -5.312253e-013, 5.124285e-011, 5.702935e-009,
  2.7652e-011, -1.093653e-012, 2.85216e-010, -2.58144e-011,
  -3.559556e-012, -1.59318e-013, -4.924823e-011, 4.710396e-009,
  2.051068e-011, 3.770161e-014, 1.311408e-010, 9.601347e-010,
  -3.052987e-012, -8.594702e-014, -2.83167e-011, 3.869278e-009,
  1.522499e-011, 1.960859e-014, 1.054377e-010, 1.53513e-009,
  -2.383354e-012, -1.441806e-013, -7.290337e-012, 3.082512e-009,
  1.134623e-011, -2.032804e-013, 1.248049e-010, 1.894534e-009,
  -1.740396e-012, -1.749606e-013, -1.67208e-011, 2.411932e-009,
  8.487226e-012, -1.330692e-013, 5.584648e-011, 2.010888e-009,
  -1.069385e-012, -1.537013e-013, -1.665115e-011, 1.851085e-009,
  6.484563e-012, 2.825036e-014, 4.266709e-011, 2.088321e-009,
  -5.208041e-013, -1.067264e-013, -1.368346e-011, 1.391269e-009,
  4.980372e-012, -1.300286e-014, -3.18619e-012, 1.977131e-009,
  3.716274e-014, -9.742453e-014, -3.194622e-011, 1.010116e-009,
  3.924811e-012, 3.333705e-014, 5.205962e-011, 1.94929e-009,
  3.264467e-013, -1.060188e-013, -2.621102e-011, 7.212878e-010,
  3.19117e-012, 3.504092e-014, 1.656603e-011, 1.779081e-009,
  6.10056e-013, -4.098291e-014, 4.578035e-012, 5.209125e-010,
  2.642378e-012, -2.420258e-014, -1.945008e-011, 1.59412e-009,
  8.136253e-013, -2.095872e-014, 6.440044e-012, 3.42592e-010,
  2.232666e-012, -2.536669e-015, -1.160622e-012, 1.49074e-009,
  9.671534e-013, 2.024186e-014, -6.564351e-012, 1.913289e-010,
  1.928802e-012, -6.072317e-015, -1.298185e-011, 1.330733e-009,
  1.053457e-012, -3.580144e-014, -2.077547e-011, 6.728202e-011,
  1.723644e-012, -1.498842e-014, -1.155156e-011, 1.183301e-009,
  1.117945e-012, -8.135747e-015, -6.357825e-012, 1.723837e-011,
  1.560286e-012, -4.846553e-015, 2.269124e-011, 1.077575e-009,
  1.124546e-012, -2.529013e-014, -1.005771e-011, -4.751494e-011,
  1.431059e-012, -3.012792e-014, 1.205837e-012, 9.27202e-010,
  1.125722e-012, 2.368069e-014, 5.773597e-012, -6.938301e-011,
  1.340111e-012, -3.094974e-014, 1.548354e-011, 8.464993e-010,
  1.082997e-012, 1.097411e-014, 8.620029e-012, -9.19091e-011,
  1.242827e-012, 5.072414e-014, -3.813893e-011, 6.969844e-010,
  1.048201e-012, 4.405746e-014, 3.990372e-012, -1.188224e-010,
  1.189272e-012, 6.270313e-014, -2.126043e-011, 6.526732e-010,
  1.001701e-012, 1.610663e-014, 6.652424e-012, -1.156064e-010,
  1.125711e-012, 3.462051e-014, -1.725951e-011, 5.770919e-010,
  9.312321e-013, 1.497081e-014, 2.407455e-011, -9.274555e-011,
  1.111997e-012, -4.998775e-014, 7.775341e-013, 5.161531e-010,
  8.831919e-013, -7.11418e-014, 1.364031e-011, -9.398148e-011,
  1.003679e-012, -6.778282e-014, 1.193915e-012, 4.325292e-010,
  8.434299e-013, -5.070572e-014, -9.110374e-012, -1.350507e-010,
  9.684046e-013, -3.26081e-014, 3.431848e-011, 4.221385e-010,
  7.539105e-013, -1.181078e-014, 3.481314e-011, -5.184243e-011,
  9.143144e-013, -1.89722e-014, -2.919573e-013, 3.371768e-010,
  6.910495e-013, 1.648267e-014, 6.015952e-011, 1.023546e-011,
  8.517453e-013, -2.176617e-013, 3.175541e-011, 3.525921e-010,
  5.80463e-013, -8.069964e-014, 2.941719e-011, -4.614836e-011,
  7.593896e-013, 2.198768e-014, 2.69121e-012, 2.755617e-010,
  6.221739e-013, 1.641841e-014, -5.769916e-011, -1.508457e-010,
  7.466222e-013, -4.688808e-014, 1.113458e-011, 3.065786e-010,
  5.783185e-013, 2.175492e-014, 1.555594e-011, -5.615471e-011,
  7.291302e-013, -7.076172e-014, -2.628609e-011, 2.013535e-010,
  5.124171e-013, 3.839199e-015, -1.443952e-011, -1.025746e-010,
  6.951543e-013, 1.695492e-014, -1.810875e-012, 2.131084e-010,
  5.367015e-013, -5.102849e-014, -3.362697e-012, -5.940535e-011,
  6.54131e-013, 4.381163e-014, 1.462329e-011, 2.119265e-010,
  4.533182e-013, -1.59816e-014, 4.328025e-012, -3.658147e-011,
  6.03179e-013, -3.263027e-014, -6.541096e-013, 1.635602e-010,
  4.075645e-013, -5.055042e-014, -1.179541e-011, -6.293114e-011,
  5.829295e-013, -3.439473e-014, 1.478586e-011, 1.737163e-010,
  3.813791e-013, -5.530276e-014, -8.523428e-012, -4.256776e-011,
  5.342047e-013, -4.1886e-014, -3.371516e-014, 1.482243e-010,
  3.592337e-013, -5.404452e-014, 2.126557e-012, -2.157836e-011,
  5.612709e-013, -4.958148e-014, 2.762668e-011, 1.614303e-010,
  3.339613e-013, -9.383132e-014, -3.264477e-011, -8.493738e-011,
  5.184769e-013, -5.253877e-014, 6.615355e-012, 1.34312e-010,
  3.06286e-013, -3.987136e-014, -2.693773e-011, -5.746434e-011,
  4.548021e-013, -7.607751e-014, -3.624179e-013, 1.258493e-010,
  3.246779e-013, -5.584655e-014, -3.795724e-011, -6.228222e-011,
  4.425811e-013, -7.714661e-014, 2.378788e-011, 1.389437e-010,
  2.737566e-013, -5.384893e-014, -5.541111e-013, -2.226986e-011,
  4.169967e-013, -4.106022e-014, 1.187967e-011, 1.152671e-010,
  2.34929e-013, 7.859415e-015, -6.969476e-012, -1.432642e-011,
  4.061129e-013, 1.196213e-014, 3.959912e-011, 1.8333e-010,
  2.706021e-013, 9.050373e-014, 1.536792e-011, 3.306675e-011,
  3.502901e-013, -2.110495e-013, -1.336338e-011, 1.011973e-010,
  1.911779e-013, -3.373771e-014, 8.0952e-012, -1.28337e-011,
  3.615553e-013, -6.942954e-014, 1.929308e-011, 1.222187e-010,
  1.792979e-013, -8.580698e-014, -2.677813e-012, -1.89155e-011,
  3.567599e-013, -6.611077e-014, 3.503464e-012, 8.938859e-011,
  3.116767e-013, -7.24954e-014, 1.689385e-011, 2.93629e-011,
  3.40178e-013, -3.018098e-014, -1.802542e-011, 5.008153e-011,
  1.98475e-013, -5.818914e-014, 2.559728e-011, 3.959346e-011,
  2.735555e-013, -9.189378e-014, -4.999189e-012, 6.586076e-011,
  1.851428e-013, -1.306308e-013, -2.646407e-011, -3.227767e-011,
  2.598907e-013, -5.813924e-014, 1.438183e-011, 8.183958e-011,
  1.556113e-013, -1.009633e-013, -1.246548e-011, -1.086856e-011,
  2.543798e-013, -1.00794e-013, 7.686295e-012, 5.221034e-011,
  1.063633e-013, -2.982328e-014, -1.635237e-012, -1.230289e-011,
  2.818109e-013, -8.471979e-014, 2.25506e-011, 7.835759e-011,
  1.43437e-013, -1.003416e-013, 4.533292e-012, -3.536124e-012,
  2.326519e-013, -1.049861e-013, 5.519001e-012, 4.407629e-011,
  1.545547e-013, -9.309928e-015, -2.169893e-011, -2.72069e-011,
  2.325462e-013, -8.235888e-014, 3.282173e-011, 9.15476e-011,
  1.632912e-013, -6.636663e-014, -1.82042e-011, -2.42848e-011,
  2.280957e-013, -4.750383e-014, 4.12585e-011, 1.089592e-010,
  8.843185e-014, -8.197046e-014, -6.89669e-012, -1.281478e-011,
  1.718178e-013, 3.008153e-015, 4.976882e-011, 1.227395e-010,
  1.185837e-013, 3.572946e-014, 2.010581e-011, 2.325531e-011,
  1.638948e-013, -2.813868e-014, 1.367619e-011, 6.370965e-011,
  1.214052e-013, -4.520589e-014, 2.768878e-012, 7.640479e-013,
  1.635846e-013, -2.742891e-014, 5.044565e-012, 4.508837e-011,
  1.205007e-013, -1.359709e-014, 1.648718e-011, 1.835521e-011,
  1.71014e-013, -4.762912e-014, 6.374493e-012, 5.350321e-011,
  1.02195e-013, 1.339422e-014, -4.902469e-012, -1.845956e-011,
  1.687618e-013, -2.498269e-014, -5.415887e-013, 3.846974e-011,
  1.102622e-013, -9.990834e-016, -6.799787e-012, -2.204746e-011,
  1.688876e-013, -1.234655e-015, 4.450934e-012, 4.54705e-011,
  1.001822e-013, -3.860124e-015, -4.89924e-012, -1.568109e-011,
  1.49982e-013, -4.818565e-014, 2.613147e-012, 4.179412e-011,
  8.588637e-014, -2.115893e-014, -2.63953e-011, -4.650782e-011,
  1.470415e-013, -6.64987e-014, -4.51778e-012, 5.034084e-011,
  7.696942e-014, -7.010123e-014, -3.026501e-011, -4.48458e-011,
  1.443204e-013, -3.378942e-014, -1.759157e-011, 1.801837e-011,
  2.563967e-014, 1.521008e-014, -3.731707e-011, -4.515188e-011,
  1.156337e-013, -1.997707e-014, -2.863603e-011, 9.247889e-012,
  7.936469e-014, -8.607242e-014, -7.35195e-012, -4.861984e-012,
  1.232301e-013, 2.592697e-014, 1.339308e-011, 6.288747e-011,
  1.355802e-013, 3.628171e-014, 4.544951e-011, 3.934498e-011,
  1.285607e-013, 1.733315e-014, 2.890037e-011, 5.633934e-011,
  1.408272e-013, -9.626939e-014, 7.462013e-011, 6.584531e-011,
  2.361384e-013, -9.878627e-014, 9.866639e-011, 1.753248e-010,
  1.158822e-013, -7.546499e-014, 1.617285e-012, 8.774134e-012,
  3.294847e-014, -6.204237e-014, 9.365776e-012, 3.465356e-011,
  1.682965e-014, -4.576838e-014, -1.400556e-011, 1.427699e-011,
  8.8668e-014, -9.009524e-014, -2.895331e-015, 4.242396e-012,
  1.482801e-014, -4.545646e-013, -1.425138e-011, 2.347287e-011,
  1.401943e-013, -2.140711e-013, 9.137281e-011, 6.603693e-011,
  4.145388e-014, 1.013649e-013, 1.40422e-011, -2.376556e-012,
  -6.380074e-015, -1.557372e-013, -1.604237e-010, -2.202509e-010,
  2.163815e-013, -4.342623e-014, 7.419569e-011, 8.644586e-011,
  3.01751e-014, -7.287382e-014, -7.446476e-011, -9.979807e-011,
  -1.373801e-014, -4.827424e-014, -9.728907e-011, -1.79866e-010,
  7.316558e-014, -5.892102e-014, -6.857426e-011, -8.354804e-011,
  2.411871e-013, -1.91542e-013, 7.229765e-011, 9.774581e-011,
  2.456728e-013, -8.901018e-015, 2.419652e-010, 3.358746e-010,
  1.065607e-013, -1.698282e-013, 5.202731e-011, 4.025628e-011,
  1.01804e-013, -9.993305e-016, 9.897884e-011, 1.685033e-010,
  1.974984e-013, -1.942199e-013, 1.4455e-010, 1.618178e-010,
  2.019318e-013, -4.308896e-014, 2.64576e-010, 3.936724e-010,
  7.482223e-015, -6.115509e-015, 1.258572e-011, 2.055776e-011,
  7.378892e-016, -1.944741e-014, 4.304835e-011, 6.43344e-011,
  4.306881e-015, -5.468029e-014, -8.61797e-011, -1.11262e-010,
  5.02187e-013, -1.96073e-013, 4.143519e-010, 5.351984e-010,
  1.663202e-013, -4.307738e-014, 1.117354e-010, 1.445906e-010,
  1.030989e-013, -7.258189e-014, 1.109109e-010, 1.446158e-010,
  1.610755e-013, -5.291206e-014, 5.964091e-011, 4.726642e-011,
  1.277972e-013, -5.033844e-014, 7.409882e-011, 1.035311e-010,
  7.918851e-014, 3.19027e-014, 3.268111e-011, 3.242622e-011,
  6.358977e-014, -1.583585e-014, 6.6296e-011, 1.074001e-010,
  4.317106e-014, -1.090365e-014, 6.691213e-012, -1.82836e-012,
  4.705004e-014, -7.26977e-014, 1.466426e-011, 6.755499e-012,
  3.453151e-014, -1.098049e-014, -1.619906e-011, -4.176515e-011,
  2.194608e-014, -2.893212e-014, 1.168454e-011, 1.69201e-011,
  7.725113e-014, -3.179575e-014, 1.038809e-011, 5.819259e-012,
  1.12841e-013, -5.27967e-014, 1.169849e-011, 2.492148e-011,
  1.406622e-013, -5.091588e-014, -1.748069e-011, -3.157122e-011,
  7.391886e-014, -2.546477e-014, -5.42549e-011, -3.989271e-011,
  5.79953e-014, -1.570965e-014, -8.628069e-012, -2.926132e-011,
  8.204444e-014, -4.329743e-014, -6.120268e-012, 1.625819e-011,
  2.021055e-014, -3.15685e-014, 7.27162e-013, -5.759815e-013,
  4.890843e-014, -1.121206e-014, 1.361502e-011, 3.099216e-011,
  4.24975e-014, -2.770784e-014, 5.944165e-012, 1.084579e-011,
  6.058539e-014, -1.555243e-014, 6.260229e-012, 1.909929e-011,
  1.013572e-013, -8.018317e-016, 2.427147e-011, 2.393838e-011,
  5.681667e-014, -4.230346e-014, -1.975653e-011, -2.855507e-011,
  6.222493e-014, -2.232883e-014, -1.495559e-011, -3.762539e-011,
  5.210129e-014, -1.744186e-014, -8.936144e-012, -5.218018e-012,
  4.282775e-014, -8.055425e-015, -8.998263e-012, -8.1917e-012,
  4.770632e-014, -2.786038e-014, -8.520847e-014, -4.155371e-012,
  3.980346e-014, 1.894912e-014, -3.877437e-011, -7.05242e-011,
  5.062745e-014, -1.460348e-014, 1.461129e-011, 2.548813e-011,
  9.636926e-014, -5.337137e-015, 2.137427e-013, -1.47922e-011,
  5.709782e-014, -3.241338e-014, 8.947306e-012, 1.150631e-011,
  7.633045e-014, -2.55167e-014, -1.235413e-011, -7.10917e-012,
  4.316645e-014, 8.332394e-015, -2.170726e-011, -3.458024e-011,
  3.933597e-014, -8.227329e-015, 1.521541e-011, 2.380597e-011,
  1.102272e-013, -4.438753e-014, 4.132302e-012, -5.878385e-013,
  6.555613e-014, 1.908032e-014, 4.119287e-011, 5.430856e-011,
  9.381143e-014, -2.494263e-014, 2.27301e-011, 7.431438e-012,
  4.728718e-014, -2.66456e-014, 8.245907e-012, 1.507635e-011,
  5.912238e-014, -4.989642e-014, -8.004262e-012, -3.039189e-012,
  3.002059e-014, 1.554154e-014, -1.988757e-011, -2.640465e-011,
  1.000265e-013, -4.897167e-014, -1.456635e-011, -1.787127e-011,
  1.126436e-013, 1.373052e-014, 3.74087e-011, 2.330888e-011,
  2.773969e-013, -9.643579e-014, 2.021863e-010, 2.783873e-010,
  9.282227e-014, -3.336821e-015, -2.628866e-011, -5.89773e-011,
  8.882856e-014, -9.014674e-014, 7.916939e-011, 1.063316e-010,
  -4.372548e-015, -3.695144e-014, -4.764507e-011, -6.306293e-011,
  2.833154e-014, -7.781124e-014, -2.014731e-011, -1.965751e-011,
  6.815545e-014, 2.503755e-014, -1.039111e-010, -1.046261e-010,
  1.541156e-013, -3.144928e-014, 2.727389e-011, 2.755472e-011,
  -2.056975e-014, 1.483217e-014, -7.787444e-011, -1.035288e-010,
  4.693905e-014, -3.783259e-014, -1.105623e-011, -1.582366e-011,
  5.7793e-014, 4.04491e-015, 7.749428e-011, 9.387203e-011,
  -5.053254e-014, -4.240863e-015, -2.359979e-011, -9.60903e-012,
  9.122978e-014, 1.887148e-014, 7.243564e-011, 7.154349e-011,
  9.022022e-014, -2.002715e-014, -5.839447e-012, -1.220671e-011,
  8.792848e-014, -1.532561e-014, 9.442021e-011, 1.095704e-010,
  -2.968926e-014, -4.636571e-014, -8.822919e-011, -1.143187e-010,
  -5.317193e-014, -1.259019e-015, -9.580379e-012, -2.668547e-011,
  -2.491514e-015, -3.528341e-014, -5.260224e-011, -5.753362e-011,
  -2.341194e-013, 7.243034e-014, -2.5251e-010, -3.473771e-010,
  -3.579368e-014, -4.160852e-014, -1.683713e-010, -2.32459e-010,
  2.442684e-013, 3.02324e-015, 1.917218e-010, 2.602721e-010,
  -1.247184e-014, 1.236142e-014, 1.991224e-011, 6.315688e-012,
  -8.214407e-014, 6.251656e-015, 1.195953e-010, 1.684487e-010,
  -6.488335e-014, -2.253223e-014, 6.66759e-011, 8.055054e-011,
  -3.933146e-014, 4.100751e-014, -3.763587e-011, -2.659896e-011,
  2.492039e-014, -7.160077e-014, -4.235548e-011, -7.662195e-011,
  2.635978e-013, 6.355838e-014, 2.345681e-010, 3.274609e-010,
  8.358074e-015, 1.863699e-014, 5.484492e-011, 7.967763e-011,
  -6.645247e-014, 8.048915e-014, -5.11153e-011, -7.81311e-011,
  -1.1794e-013, -7.037648e-014, -1.070452e-010, -1.125372e-010,
  -5.776255e-013, 1.060414e-013, -6.633424e-010, -9.242731e-010,
  1.803793e-013, -9.034371e-014, 1.401932e-010, 2.62546e-010,
  -7.214153e-014, -1.526388e-014, -1.281917e-010, -1.869503e-010,
  1.465825e-013, -8.138969e-014, 9.417533e-011, 1.118692e-010,
  1.201114e-014, -1.70773e-015, -1.589688e-011, -3.62566e-011,
  2.402986e-014, -4.744989e-014, -5.380183e-011, -6.828874e-011,
  -1.017649e-014, -3.837482e-016, -2.733034e-011, -1.046718e-011,
  7.849855e-014, 1.316632e-016, -2.358165e-011, -3.5573e-011,
  1.354771e-013, 3.202232e-014, 5.852899e-011, 6.466462e-011,
  7.025499e-014, 1.986358e-014, 3.380521e-011, 4.707013e-011,
  3.469409e-014, -2.674294e-014, -2.129965e-011, -2.597273e-011,
  8.498871e-014, -1.813869e-014, -1.295703e-011, -2.488002e-011,
  4.727117e-014, -3.383118e-014, -1.772699e-011, -3.373905e-011,
  2.671429e-014, -6.818423e-015, 2.121984e-011, 3.546959e-011,
  3.634862e-014, 3.122161e-014, 1.731073e-011, 2.750678e-011,
  -1.08804e-015, -4.641107e-014, -4.687778e-013, -7.983676e-012,
  2.618301e-014, 2.291837e-014, 2.723713e-011, 3.810875e-011,
  -3.575434e-014, -2.299359e-014, -6.604826e-012, -1.572824e-011,
  -7.542483e-014, -4.76093e-015, 3.180275e-012, -1.377487e-011,
  7.479409e-014, -2.802438e-014, -5.395706e-012, -1.102164e-011,
  -2.184645e-014, -1.49159e-014, 8.189049e-012, 1.779862e-012,
  -2.190487e-014, -2.703281e-014, -2.402301e-011, -3.681539e-011,
  1.127426e-013, -1.008147e-014, 8.927213e-011, 1.376667e-010,
  5.416986e-014, 5.181486e-014, 7.230261e-011, 1.107375e-010,
  1.874394e-013, -5.409271e-015, 3.707334e-011, 1.024423e-010,
  1.072702e-013, 1.147857e-016, 1.55097e-010, 1.896267e-010,
  7.380111e-015, -3.988041e-014, -4.240963e-011, -9.072036e-011,
  6.9601e-014, -5.989186e-014, 9.299316e-012, 1.642344e-012,
  7.064791e-014, -3.219004e-014, 5.592492e-011, 5.955589e-011,
  1.14297e-015, 2.651063e-015, 4.721936e-011, 6.754799e-011,
  5.346371e-014, -4.646007e-014, 2.186231e-012, 3.643657e-011,
  -4.983786e-014, -6.8422e-014, 3.026621e-011, 4.552928e-011,
  -1.307683e-013, -5.682413e-014, -6.610693e-011, -7.261135e-011,
  -9.852704e-014, 3.819019e-014, -8.179824e-011, -1.339696e-010,
  -5.183218e-014, -5.27307e-015, -1.127072e-010, -1.383464e-010,
  -3.333381e-014, -4.045689e-014, -1.04749e-011, 1.270503e-011,
  5.395325e-014, -7.177032e-014, -3.220658e-011, -3.08694e-011,
  1.836231e-013, -6.361381e-014, 1.579284e-010, 2.150461e-010,
  -2.862934e-014, 1.547853e-014, -1.379945e-011, -1.880252e-011,
  1.970037e-014, 1.715408e-015, -5.023248e-011, -6.618164e-011,
  3.670178e-014, -2.231794e-014, -2.348587e-011, -4.157288e-012,
  1.290504e-013, 2.738477e-014, 7.791134e-011, 9.586232e-011,
  -8.068252e-015, -2.102498e-014, -4.053147e-012, 6.697974e-012,
  -4.35689e-014, 1.135527e-014, 4.418387e-011, 5.917918e-011,
  -1.045496e-013, 1.00801e-013, -1.868962e-011, -1.844666e-011,
  -7.66899e-014, -8.475056e-014, 6.709626e-011, 5.757346e-011,
  6.332428e-015, 4.932087e-014, 5.756982e-012, -5.436047e-012,
  1.068076e-013, -3.886171e-014, 5.417904e-012, 2.69455e-012,
  4.483142e-014, -2.868102e-014, 3.336729e-011, 3.921774e-011,
  9.477038e-014, -5.224526e-014, 2.830834e-011, 4.072018e-011,
  -1.351158e-014, 1.746756e-014, -3.04446e-011, -3.026059e-011,
  -8.339304e-015, 6.964151e-014, 3.003528e-011, 4.139934e-011,
  6.318107e-014, 1.097397e-014, 1.586717e-011, 3.559013e-011,
  -3.312183e-014, -2.468487e-014, 3.004834e-011, 3.910688e-011,
  -2.554082e-014, -1.752923e-015, -5.578809e-011, -8.88311e-011,
  -3.69718e-014, -2.625016e-014, -3.460069e-011, -4.880322e-011,
  -6.841159e-015, -6.463912e-015, 3.129057e-011, 3.990239e-011,
  2.304735e-014, 1.022053e-016, 1.326548e-012, -5.785406e-012,
  -4.312117e-014, -3.642412e-014, -4.437642e-011, -5.688982e-011,
  -4.261101e-014, -7.576824e-016, 1.188495e-011, 4.343571e-011,
  -6.721181e-014, -8.767796e-015, -4.261722e-013, 1.406548e-012,
  -2.089075e-014, -2.481146e-014, 6.092426e-012, 3.653483e-011,
  -1.500112e-014, -6.329584e-015, -5.15625e-012, -1.118471e-011,
  -9.079693e-016, 2.506391e-014, 4.420991e-012, 1.694521e-011,
  2.610909e-014, 5.484457e-014, 2.458653e-011, 1.293005e-011,
  4.856781e-014, 2.936155e-014, -3.064726e-011, -4.813328e-011,
  5.598144e-014, 4.161566e-015, 3.82364e-011, 7.160225e-011,
  7.893314e-016, 4.001172e-015, 1.892656e-012, -4.96823e-012,
  8.398865e-015, 2.579716e-014, -3.204016e-011, -1.207247e-011,
  3.365585e-014, -3.356474e-014, 1.250596e-010, 1.484888e-010,
  6.56613e-014, -5.629102e-014, 8.772294e-011, 1.339719e-010,
  -1.703534e-014, 4.692464e-014, -1.628552e-011, -1.631818e-011,
  3.456506e-013, -5.338472e-014, 3.448515e-010, 4.301569e-010,
  8.73348e-014, 6.757331e-014, 1.28697e-010, 2.006384e-010,
  1.623797e-013, 2.90295e-014, 9.4215e-011, 1.507077e-010,
  2.805232e-013, 3.245741e-014, 4.429309e-010, 6.311821e-010,
  -1.430424e-014, -3.595964e-014, -8.330373e-011, -1.278674e-010,
  3.627673e-014, -4.093323e-014, 9.667576e-011, 1.429477e-010,
  1.918299e-013, -2.387396e-014, 3.471912e-010, 4.649648e-010,
  -1.975567e-013, -3.654737e-015, -8.215337e-011, -1.253745e-010,
  -7.04981e-014, 1.963282e-014, -1.508864e-010, -2.308522e-010,
  -2.081148e-013, 2.809621e-014, -3.589983e-010, -4.77182e-010,
  -1.238658e-013, -2.202686e-014, -2.462458e-010, -3.521139e-010,
  1.690774e-013, -1.323451e-014, 2.812699e-011, 5.366269e-011,
  -9.553273e-014, 6.339563e-014, -7.356643e-011, -9.804162e-011,
  -8.021856e-015, -2.94448e-014, -8.828743e-011, -1.403214e-010,
  -9.484445e-014, 3.44011e-014, -1.005981e-010, -1.329204e-010,
  2.28735e-014, -7.10974e-014, -4.394405e-011, -6.106943e-011,
  -7.868292e-014, 2.8109e-014, -2.019743e-011, -1.68929e-011,
  -1.045542e-013, 7.305549e-014, -1.140165e-010, -1.854645e-010,
  -4.438574e-014, -1.508099e-015, -2.280028e-011, -1.840267e-011,
  4.060666e-014, -2.505777e-014, 3.614848e-012, 1.367924e-011,
  1.010401e-015, 7.952945e-014, -2.110876e-011, -4.161162e-011,
  1.259888e-013, -4.974552e-015, 7.922421e-012, 3.156754e-011,
  1.344132e-013, 4.554675e-014, 1.108986e-010, 1.433191e-010,
  5.102476e-014, 1.774606e-015, 1.187709e-010, 1.576506e-010,
  -6.953803e-015, -2.566834e-014, -4.897961e-011, -5.934048e-011,
  1.37446e-013, -2.014821e-014, 8.15724e-011, 1.087135e-010,
  -1.13036e-013, 4.778864e-014, -9.248417e-011, -1.249948e-010,
  -4.191684e-014, -2.305873e-014, -8.330242e-012, -5.304352e-012,
  -2.72049e-014, -2.416867e-014, -4.473604e-011, -5.241694e-011,
  5.046411e-014, -5.409029e-014, -3.485169e-011, -1.31683e-011,
  2.612223e-014, -6.723713e-014, -4.243452e-011, -9.81601e-011,
  8.857766e-014, -4.993655e-014, 7.812283e-011, 1.02659e-010,
  1.913427e-014, 3.535352e-014, -4.038812e-011, -4.384867e-011,
  -6.990495e-014, -1.707597e-014, -2.295359e-011, -4.516543e-011,
  1.301769e-014, -1.561885e-015, 3.303386e-011, 7.230267e-011,
  -2.290749e-014, -6.689277e-014, -1.503156e-011, -5.755008e-012,
  5.940603e-014, -1.743277e-014, 2.567807e-011, 4.65145e-011,
  -6.407584e-014, 3.609296e-015, -1.1509e-010, -1.320346e-010,
  -2.610921e-014, -2.826828e-014, -1.644731e-011, -2.915434e-011,
  -8.253324e-014, 5.920846e-014, -4.79866e-011, -5.296287e-011,
  -2.02862e-013, 7.989622e-015, -2.548287e-010, -3.441784e-010,
  -1.273194e-014, 2.553601e-014, -6.201793e-011, -1.110316e-010,
  2.381924e-013, -3.399777e-014, 3.265082e-010, 4.707104e-010,
  2.078718e-014, -1.243097e-014, 1.695293e-010, 2.285026e-010,
  2.650552e-013, -8.390032e-014, 1.958684e-010, 3.011217e-010,
  4.031539e-014, 1.258685e-014, 2.960504e-010, 3.419539e-010,
  1.341958e-013, -5.491997e-014, 5.068379e-011, 7.923354e-011,
  3.38206e-013, 5.836964e-014, 5.613577e-010, 7.537709e-010,
  1.35294e-013, -3.740286e-014, 7.545288e-011, 1.407626e-010,
  -4.153927e-014, 5.394007e-014, 3.016755e-011, 5.037601e-011,
  -1.609691e-014, 1.010364e-013, 1.271125e-010, 1.298607e-010,
  -5.013227e-013, 1.623923e-013, -6.962192e-010, -9.581624e-010,
  -5.026236e-013, 5.095508e-014, -7.26752e-010, -9.346247e-010,
  3.35268e-013, -9.793068e-014, 5.153789e-010, 7.431848e-010,
  -4.905385e-013, 3.648337e-014, -6.591788e-010, -8.879475e-010,
  2.123363e-013, -9.965353e-014, 2.572769e-010, 4.055433e-010,
  1.899335e-014, 5.821273e-016, 6.928929e-014, -2.256952e-012,
  1.922979e-014, 3.62264e-016, -3.622752e-012, 2.12796e-012,
  1.851101e-015, 3.800039e-015, 2.763519e-011, 1.85122e-011,
  5.357106e-015, 2.504035e-015, 7.234197e-012, 1.610133e-011,
  -4.877318e-014, 1.042475e-014, -3.258505e-012, -2.094768e-012,
  -2.634775e-014, 6.671186e-015, 9.939269e-012, 1.316271e-011,
  3.949384e-015, 5.838382e-016, -1.89074e-011, -2.752509e-011,
  1.61591e-014, -1.702493e-014, -6.863459e-012, 4.407648e-012,
  2.338566e-014, -2.150998e-015, -2.026748e-012, -4.35034e-012,
  2.31492e-014, 3.645353e-015, 1.277903e-012, 7.140041e-012,
  2.161098e-014, 7.11855e-016, 7.201593e-012, 1.465878e-011,
  2.520007e-014, 1.324143e-015, 1.909082e-012, 1.086303e-011,
  5.276429e-014, -1.110526e-014, 5.569376e-012, 2.421157e-012,
  -5.030095e-014, 1.458757e-014, 7.094168e-013, 7.882648e-012,
  1.132229e-014, -1.904452e-014, -9.807011e-012, -1.78386e-011,
  2.080666e-014, -6.10252e-015, 7.021044e-012, 1.87847e-011,
  3.561815e-014, -1.794402e-015, 4.683702e-011, 3.651704e-011,
  4.419444e-014, 5.767064e-016, 3.082321e-012, 1.374537e-011,
  5.664514e-014, 1.364271e-013, 4.446098e-011, 3.640782e-011,
  5.375378e-014, 9.012349e-014, 3.549048e-012, 1.524888e-011,
  3.928047e-014, 3.551258e-015, 9.17766e-012, 1.101966e-011,
  1.114246e-013, -9.048918e-015, -7.280821e-012, 3.316262e-013,
  3.073873e-014, -1.635902e-016, -6.557356e-013, -1.372526e-012,
  3.370508e-014, 6.718795e-016, -1.205513e-012, 5.977172e-012,
  3.050142e-014, 2.017947e-016, 7.836257e-012, 4.049025e-012,
  2.854084e-014, -1.38911e-016, 4.446618e-012, 1.195299e-011,
  2.799026e-014, -2.120762e-015, -1.728986e-012, -5.177078e-012,
  2.392704e-014, 3.296155e-015, -1.139875e-011, -2.686315e-012,
  3.161203e-014, -5.631483e-016, -3.786325e-012, -6.438962e-012,
  2.564717e-014, 2.573217e-015, -5.987293e-012, 2.114762e-012,
  2.00215e-014, 2.868269e-015, 7.094188e-012, 8.874653e-012,
  3.63571e-014, 2.993237e-015, 3.393195e-012, 1.669729e-011,
  7.506821e-014, -3.691525e-015, 6.112633e-011, 8.119149e-011,
  6.493643e-014, 4.611515e-015, -2.266074e-011, -1.59054e-011,
  2.616912e-014, 3.131347e-015, -3.227432e-012, -6.040697e-012,
  3.139115e-014, 5.72768e-015, -3.164726e-013, 1.187475e-011,
  2.677187e-014, 1.872751e-014, -2.842197e-012, -6.52464e-012,
  3.026305e-014, -2.302345e-015, 2.28403e-013, 1.146544e-011,
  3.258082e-014, 9.598482e-015, 1.045358e-011, 1.14308e-011,
  3.687204e-014, -1.921166e-015, -7.933894e-012, 3.975747e-012,
  3.979239e-014, -1.477746e-015, 2.469906e-011, 2.898879e-011,
  4.972607e-014, 1.976079e-015, -1.106785e-011, 3.649142e-012,
  2.464469e-014, 1.482116e-017, 8.565925e-012, 5.841693e-012,
  4.576293e-014, -2.568082e-015, -1.698306e-012, 1.136279e-011,
  2.323514e-014, 1.640982e-015, -3.059561e-011, -4.287387e-011,
  1.074672e-014, 2.913654e-015, -1.323338e-012, 1.404253e-011,
  7.007322e-014, -1.075492e-014, -1.824303e-011, -2.360382e-011,
  3.429211e-014, -3.188682e-015, 1.325236e-012, 1.806507e-011,
  2.990928e-014, -5.04228e-015, -5.36264e-013, 4.517573e-012,
  4.247985e-014, -4.293328e-015, 6.7008e-012, 2.221373e-011,
  2.778456e-014, -3.772067e-015, -8.333134e-012, -9.877441e-012,
  3.981461e-014, -3.097824e-015, 2.695291e-012, 1.238867e-011,
  3.981057e-014, -8.208719e-015, -9.974139e-012, -1.37532e-011,
  4.532286e-014, 1.013673e-015, -6.792059e-012, 4.688758e-012,
  -5.772504e-014, 1.092566e-014, -4.96608e-012, -5.785833e-012,
  1.75826e-014, 2.671559e-015, 2.46705e-011, 2.884666e-011,
  2.116647e-014, -3.274227e-016, 7.634318e-013, 4.485295e-012,
  4.795569e-014, 3.215443e-015, 8.014937e-012, 1.945857e-011,
  2.026134e-014, -1.242399e-015, 2.525542e-011, 2.857086e-011,
  7.235465e-014, -3.263578e-015, 2.085447e-011, 3.708392e-011,
  3.495242e-014, -3.319209e-015, 1.706851e-012, -5.181969e-012,
  4.821242e-014, -4.209107e-015, 4.088088e-013, 1.371279e-011,
  4.871865e-014, -2.329764e-015, -8.115595e-012, 5.084101e-012,
  5.122808e-014, -7.21392e-015, -5.501814e-012, 2.552523e-011,
  4.723222e-014, -2.252593e-015, 2.095015e-012, 1.273682e-012,
  5.191437e-014, -3.895717e-015, -1.26678e-012, 1.197511e-011,
  1.773862e-014, 1.770302e-015, 2.407217e-012, 8.122138e-012,
  3.791646e-014, -2.96557e-015, 3.306104e-012, 1.858899e-011,
  3.511339e-014, -1.913881e-015, -4.090367e-013, 1.804142e-012,
  5.119642e-014, -1.306898e-015, -7.403069e-012, 1.035806e-011,
  -2.127644e-016, -1.827812e-015, -4.960562e-012, -1.315537e-011,
  -2.035344e-015, -1.767163e-015, 4.484214e-012, 1.860515e-011,
  -6.059929e-015, 2.536667e-015, -3.168485e-011, -4.661972e-011,
  -2.871032e-014, 2.879789e-015, 7.774725e-013, 1.694332e-011,
  3.853008e-014, -8.959795e-016, 2.889455e-012, -4.38101e-013,
  6.673008e-014, -7.115302e-015, 1.004612e-011, 2.808888e-011,
  3.407021e-014, -2.766598e-015, -1.295828e-012, -6.277275e-012,
  6.155454e-014, -6.65512e-015, -1.365568e-012, 1.504168e-011,
  4.678066e-014, -5.00041e-015, -2.722922e-014, -4.528197e-012,
  8.105139e-014, -4.538047e-015, -1.823074e-012, 1.701005e-011,
  9.239376e-014, -6.768392e-015, 3.747498e-012, -3.22484e-012,
  1.252182e-013, -7.929069e-015, -2.410259e-013, 2.031825e-011,
  6.198697e-014, -3.539276e-015, 2.132466e-011, 1.952819e-011,
  8.821986e-014, 1.32035e-015, 4.790157e-012, 3.385945e-011,
  4.85101e-014, -1.75866e-015, 4.657442e-012, 1.262686e-012,
  7.665726e-014, -1.087989e-015, -3.084224e-012, 1.757139e-011,
  5.115366e-014, 1.957335e-016, -1.004754e-012, -5.669562e-012,
  7.433129e-014, 3.891241e-015, 1.412067e-014, 2.406467e-011,
  -3.016299e-014, 1.747209e-014, 1.970563e-012, -3.026598e-012,
  3.84927e-014, 1.395747e-014, 1.57295e-012, 2.704345e-011,
  4.75604e-014, 2.136169e-015, 1.352142e-012, -2.042632e-012,
  7.675613e-014, 2.669993e-015, 3.295022e-012, 2.255546e-011,
  5.929007e-014, 2.166261e-014, 4.447061e-012, -3.201405e-012,
  7.929227e-014, 2.62481e-016, -6.998049e-012, 1.330547e-011,
  5.795845e-014, 9.487134e-015, -1.458273e-012, -7.809696e-012,
  8.095284e-014, 1.312736e-014, -7.845313e-012, 1.952249e-011,
  -4.397032e-014, 4.192851e-014, 1.085783e-011, 1.230956e-011,
  1.614048e-013, 2.688602e-014, 6.358822e-012, 4.919952e-011,
  4.6609e-014, 1.373911e-014, -5.881967e-012, -3.39791e-012,
  1.045116e-013, 1.723805e-014, 2.530609e-011, 5.641772e-011,
  6.451575e-014, 1.727091e-014, -1.748672e-012, -6.807841e-012,
  9.605951e-014, 1.282881e-014, -2.767677e-012, 2.816931e-011,
  6.533969e-014, 9.031313e-015, 2.369915e-012, -5.027159e-012,
  9.560738e-014, 1.279143e-014, -7.152175e-012, 2.672263e-011,
  3.765503e-014, 1.345635e-014, 1.501631e-012, -7.56463e-012,
  7.214481e-014, 1.565537e-014, -9.190715e-012, 2.701724e-011,
  5.243312e-014, 1.734356e-014, -3.497904e-012, -1.085921e-011,
  8.465787e-014, 1.746426e-014, -7.252954e-012, 2.990858e-011,
  8.289873e-014, 1.005268e-014, -9.281032e-014, -5.813273e-012,
  1.085279e-013, 8.047237e-015, -4.965417e-012, 3.191905e-011,
  8.004951e-014, 3.68202e-015, -3.420211e-012, -1.152459e-011,
  1.094816e-013, 8.382024e-015, -9.313693e-012, 2.420697e-011,
  9.392418e-014, -2.284774e-015, 3.934385e-013, -7.776842e-012,
  1.237165e-013, 5.985416e-015, 2.13208e-012, 3.833067e-011,
  1.42248e-013, -6.013524e-015, -4.583369e-012, -1.369942e-011,
  1.257518e-013, 7.707839e-015, -3.593152e-012, 3.217083e-011,
  9.334427e-014, 3.690512e-015, 1.022115e-012, -6.555252e-012,
  1.302907e-013, 1.339433e-015, -1.407261e-012, 3.749959e-011,
  9.765446e-014, -1.138051e-015, -1.882262e-012, -7.841955e-012,
  1.364008e-013, -2.445782e-015, 9.043355e-013, 4.225252e-011,
  9.501874e-014, -2.864328e-015, -2.914446e-012, -7.812377e-012,
  1.3866e-013, -4.249242e-015, -8.896286e-013, 4.062486e-011,
  1.017119e-013, -5.460044e-015, -2.357002e-012, -8.168913e-012,
  1.462533e-013, -6.703873e-015, 6.149861e-012, 4.665398e-011,
  1.073037e-013, -4.610186e-015, 1.776432e-012, -8.050679e-012,
  1.576879e-013, -7.556275e-015, 2.726535e-012, 4.866458e-011,
  1.120651e-013, -2.343373e-015, -3.938136e-013, -8.039798e-012,
  1.587332e-013, -6.855484e-015, -1.652846e-012, 4.734194e-011,
  1.153013e-013, -3.158191e-015, -1.682956e-012, -1.046496e-011,
  1.688267e-013, -1.080324e-014, 4.055601e-012, 5.234752e-011,
  1.331771e-014, 7.091552e-015, -7.884353e-013, -6.40584e-012,
  2.265367e-013, -1.568161e-014, -1.085937e-012, 4.70478e-011,
  1.231533e-013, -1.406189e-015, -3.328698e-012, -8.413358e-012,
  1.81458e-013, -6.746269e-015, -1.382082e-012, 5.194862e-011,
  1.336288e-013, 4.472833e-016, -7.49335e-012, -1.563068e-011,
  1.912915e-013, -1.832118e-014, -2.512542e-013, 5.629496e-011,
  1.455569e-013, 2.445397e-015, -1.106795e-012, -8.83412e-012,
  2.035839e-013, -8.525868e-015, -1.766455e-012, 6.102008e-011,
  2.206475e-013, -1.711655e-014, 3.103018e-012, -6.078975e-012,
  1.724962e-013, 5.772666e-015, 5.832061e-012, 7.102454e-011,
  1.730559e-013, -9.934301e-015, -1.349791e-013, -1.174772e-011,
  2.071235e-013, -6.898355e-015, -8.351928e-013, 5.955812e-011,
  1.695299e-013, -6.464118e-015, -3.134318e-011, -3.557333e-011,
  2.311746e-013, -1.04891e-014, 6.702697e-012, 7.091647e-011,
  1.745805e-013, -7.603091e-015, -4.52564e-012, -2.019068e-011,
  2.440953e-013, -9.860252e-015, 4.854128e-012, 7.218517e-011,
  2.184801e-013, -8.495172e-015, 1.196397e-012, -1.198756e-011,
  2.772092e-013, -1.718502e-014, 4.298031e-012, 8.041057e-011,
  2.418665e-013, -1.581878e-014, 2.768523e-013, -1.306189e-011,
  2.860383e-013, -1.377579e-014, 4.243738e-012, 8.603071e-011,
  1.99908e-013, -3.818242e-015, 1.786351e-012, -1.236325e-011,
  2.965856e-013, -5.286862e-015, 3.701548e-012, 9.094395e-011,
  2.120761e-013, 5.359058e-016, 1.668477e-012, -1.349864e-011,
  3.131691e-013, -6.63768e-017, 8.698433e-014, 9.288964e-011,
  2.351406e-013, -1.261265e-015, -5.404086e-012, -2.318187e-011,
  3.213768e-013, -7.367953e-015, -1.635204e-011, 7.853564e-011,
  2.403184e-013, -4.819647e-015, -1.113258e-011, -2.954833e-011,
  3.36859e-013, -9.103369e-015, -2.093971e-011, 7.114322e-011,
  2.430603e-013, -5.74172e-015, -1.37682e-011, -2.978622e-011,
  3.783537e-013, -2.451569e-014, 9.501548e-012, 1.164547e-010,
  2.748164e-013, -5.024655e-015, -2.14478e-011, -4.162855e-011,
  3.889498e-013, -1.728448e-014, -1.949643e-012, 1.061547e-010,
  2.788682e-013, -3.549774e-015, 2.428521e-011, 1.258572e-011,
  4.424206e-013, -1.111285e-014, 1.726263e-011, 1.393691e-010,
  1.654599e-013, 2.32107e-014, -1.554603e-011, -4.429464e-011,
  4.771618e-013, -1.817637e-014, 1.715477e-011, 1.431301e-010,
  3.213083e-013, -2.040851e-015, -9.208895e-012, -3.652201e-011,
  4.640606e-013, 4.522911e-015, -2.598364e-012, 1.311769e-010,
  3.326717e-013, -4.70929e-016, -2.26557e-011, -4.898893e-011,
  5.038436e-013, -1.546926e-014, 8.690823e-012, 1.587979e-010,
  3.661487e-013, -1.094647e-014, -9.832324e-012, -3.658774e-011,
  5.418834e-013, -2.112818e-014, 1.912174e-011, 1.696155e-010,
  4.614368e-013, -2.389743e-014, 6.236963e-012, -2.454983e-011,
  5.777366e-013, -1.925604e-014, 1.120638e-011, 1.677087e-010,
  4.480158e-013, -2.303509e-014, 1.953336e-011, -9.326042e-012,
  6.577972e-013, -2.872956e-014, -6.560984e-012, 1.60798e-010,
  4.622576e-013, -2.215511e-014, -1.405687e-011, -4.906744e-011,
  6.793292e-013, -3.984175e-014, 4.50487e-012, 1.897483e-010,
  5.153889e-013, -1.437209e-014, 4.005909e-012, -3.650043e-011,
  7.452933e-013, -2.396432e-014, -6.435576e-012, 1.822398e-010,
  5.21177e-013, -3.804201e-014, -4.879415e-012, -4.853117e-011,
  8.290019e-013, -6.506236e-014, 6.465469e-012, 2.067482e-010,
  5.889291e-013, -3.608107e-014, 5.129622e-012, -5.072525e-011,
  8.924548e-013, -5.041368e-014, 5.242562e-012, 2.369091e-010,
  6.674755e-013, -2.29558e-014, 1.02077e-011, -5.026942e-011,
  9.357813e-013, -1.084386e-014, 2.068677e-011, 2.712037e-010,
  7.332161e-013, -2.695796e-015, -1.921452e-011, -9.370454e-011,
  9.895159e-013, -1.449881e-014, -4.606188e-012, 2.782667e-010,
  8.007281e-013, -3.471598e-014, 6.898366e-012, -8.612761e-011,
  1.05248e-012, -2.146113e-014, 1.23213e-011, 3.225568e-010,
  8.759569e-013, -3.433034e-014, 2.53993e-012, -1.059642e-010,
  1.136643e-012, -4.373147e-014, 1.140387e-011, 3.559848e-010,
  9.734775e-013, -2.794745e-014, 2.530087e-012, -1.270258e-010,
  1.205515e-012, -4.112704e-014, -8.696181e-013, 3.898646e-010,
  1.058432e-012, -1.953135e-014, -9.068801e-013, -1.496611e-010,
  1.276254e-012, -2.918905e-014, -7.95872e-013, 4.504404e-010,
  1.153671e-012, -1.20143e-014, -5.337356e-012, -1.643144e-010,
  1.352057e-012, -2.252107e-014, 1.890164e-012, 5.220065e-010,
  1.24464e-012, -1.886079e-014, -2.99887e-012, -1.728037e-010,
  1.442073e-012, -2.575828e-014, 6.259321e-012, 5.989422e-010,
  1.336894e-012, -8.574715e-015, 4.875782e-013, -1.764986e-010,
  1.527437e-012, 1.432034e-015, 6.651522e-013, 6.966388e-010,
  1.415913e-012, -1.845991e-014, 4.640155e-012, -1.734447e-010,
  1.618094e-012, 2.699964e-014, -6.232253e-012, 8.088377e-010,
  1.401845e-012, 2.143657e-014, 3.638722e-011, -1.186065e-010,
  1.791489e-012, 1.851711e-014, -2.385586e-011, 9.329865e-010,
  1.441688e-012, 1.316319e-014, 2.847036e-012, -1.222549e-010,
  1.870256e-012, 6.256576e-015, 4.795563e-013, 1.133642e-009,
  1.563983e-012, -6.662854e-015, 6.130554e-011, -8.73854e-012,
  1.989643e-012, 2.834798e-014, 1.029827e-011, 1.251799e-009,
  1.717513e-012, -3.224386e-014, -4.587564e-012, 2.333273e-011,
  2.1768e-012, 3.606519e-014, -1.516223e-010, 1.241748e-009,
  1.313218e-012, -2.386791e-015, 8.601763e-012, 1.819383e-010,
  2.507005e-012, 1.622863e-014, 1.264061e-011, 1.683188e-009,
  1.083349e-012, -1.420262e-014, 3.895194e-012, 3.767863e-010,
  2.926631e-012, -3.619008e-014, 2.052697e-011, 1.901107e-009,
  8.054345e-013, -3.775098e-014, 6.556279e-011, 7.243863e-010,
  3.579756e-012, -1.112157e-013, -8.404618e-012, 2.066756e-009,
  2.388965e-013, -2.647849e-014, 1.504323e-011, 1.022469e-009,
  4.462953e-012, -1.238075e-013, 4.58446e-011, 2.361714e-009,
  -4.198414e-013, -1.762441e-014, 1.193615e-011, 1.499526e-009,
  5.770222e-012, -1.472693e-013, 4.303399e-011, 2.551441e-009,
  -1.218745e-012, -1.47468e-014, 3.24183e-011, 2.1379e-009,
  7.691876e-012, -2.63997e-013, 8.136069e-011, 2.701986e-009,
  -2.187462e-012, -2.120566e-014, 5.549006e-011, 2.935465e-009,
  1.048184e-011, -4.96396e-013, 1.202978e-010, 2.707667e-009,
  -3.231396e-012, -5.181913e-014, 8.434197e-011, 3.90201e-009,
  1.447367e-011, -7.875868e-013, 1.583958e-010, 2.51987e-009,
  -4.315882e-012, -1.310428e-013, 1.21922e-010, 5.042763e-009,
  2.023455e-011, -1.23133e-012, 1.779912e-010, 1.996493e-009,
  -5.119338e-012, -2.867587e-013, 1.694752e-010, 6.411596e-009,
  2.838543e-011, -1.74199e-012, 1.474782e-010, 1.008911e-009,
  -5.045837e-012, -6.703255e-013, 2.368682e-010, 7.884961e-009,
  3.991697e-011, -2.869713e-012, 2.709536e-010, -5.035781e-010,
  -3.297435e-012, -1.396952e-012, 3.365343e-010, 9.409125e-009,
  5.614728e-011, -4.393852e-012, 3.274214e-010, -2.98844e-009,
  2.788592e-012, -2.336713e-012, 3.554055e-010, 1.079603e-008,
  7.847538e-011, -5.461933e-012, 2.717483e-010, -6.770852e-009,
  1.423084e-011, -4.204419e-012, 3.796783e-010, 1.166361e-008,
  1.114499e-010, -7.212664e-012, 2.307692e-010, -1.244078e-008,
  3.65354e-011, -7.634553e-012, 4.339789e-010, 1.129514e-008,
  1.573264e-010, -1.035465e-011, 2.566461e-010, -2.087009e-008,
  7.881121e-011, -1.197753e-011, 4.183543e-010, 8.400739e-009,
  2.233137e-010, -1.282529e-011, 2.482642e-010, -3.321494e-008,
  1.574299e-010, -1.79683e-011, 3.156962e-010, 6.43011e-010,
  3.177901e-010, -1.478884e-011, 2.501969e-010, -5.095517e-008,
  3.056484e-010, -2.596437e-011, 2.090612e-010, -1.683322e-008,
  4.566481e-010, -1.577049e-011, 4.017387e-010, -7.716141e-008,
  5.911073e-010, -3.725233e-011, 3.116108e-010, -5.337961e-008,
  6.629571e-010, -1.423534e-011, 1.049615e-009, -1.157013e-007,
  1.161002e-009, -6.727756e-011, 1.815415e-009, -1.323118e-007,
  9.700738e-010, -1.207312e-011, 3.386928e-009, -1.744527e-007,
  2.250431e-009, -1.341717e-010, 7.618936e-009, -3.138728e-007,
  1.413002e-009, -7.017024e-012, 8.281502e-009, -2.671216e-007,
  3.275153e-009, -3.095267e-010, 2.857006e-008, -7.804033e-007,
  1.843508e-009, 3.855989e-012, 1.832986e-008, -4.209459e-007,
  -2.012046e-009, -6.329687e-010, 9.2082e-008, -1.926073e-006,
  1.623923e-009, 1.972105e-011, 3.532531e-008, -6.594325e-007,
  -1.194802e-008, -6.670239e-010, 1.515176e-007, -3.294221e-006,
  1.55687e-009, 4.533373e-011, 4.300905e-008, -8.551123e-007,
  -1.398993e-008, -6.470378e-010, 1.534307e-007, -3.701134e-006,
  1.641069e-009, 1.654033e-011, 3.63718e-008, -8.983426e-007,
  -1.094965e-008, -1.051288e-009, 1.032126e-007, -3.094365e-006,
  1.92409e-009, -7.409179e-011, 2.3701e-008, -7.685331e-007,
  -5.77234e-010, -1.124077e-009, 4.024014e-008, -1.703143e-006,
  2.279222e-009, -7.056034e-011, 1.396552e-008, -5.341212e-007,
  3.370348e-009, -4.594014e-010, 1.222229e-008, -6.854856e-007,
  1.797141e-009, -2.374841e-011, 8.083029e-009, -3.568832e-007,
  2.135465e-009, -1.02756e-010, 3.408611e-009, -2.817796e-007,
  1.285058e-009, -1.635935e-012, 3.514323e-009, -2.381568e-007,
  1.096938e-009, -1.888267e-011, 6.306481e-010, -1.215977e-007,
  8.880163e-010, -2.079802e-012, 1.074471e-009, -1.599883e-007,
  5.639402e-010, -1.827298e-011, 2.205225e-010, -4.991271e-008,
  6.128675e-010, -8.958302e-012, 3.729358e-010, -1.079813e-007,
  2.959673e-010, -1.966259e-011, 3.127087e-010, -1.610984e-008,
  4.28227e-010, -1.508361e-011, 1.544151e-010, -7.325146e-008,
  1.562591e-010, -2.093093e-011, 4.999242e-010, -5.109725e-011,
  3.030608e-010, -1.832611e-011, 4.024189e-010, -4.943614e-008,
  8.000028e-011, -1.47653e-011, 6.004831e-010, 7.390768e-009,
  2.157042e-010, -1.571637e-011, 5.053782e-010, -3.297851e-008,
  3.875739e-011, -8.194192e-012, 4.411172e-010, 1.024843e-008,
  1.546275e-010, -1.03218e-011, 5.408343e-010, -2.148558e-008,
  1.634884e-011, -3.686221e-012, 3.232054e-010, 1.094237e-008,
  1.113401e-010, -5.665701e-012, 4.883695e-010, -1.346925e-008,
  4.469951e-012, -2.29066e-012, 2.98859e-010, 1.035866e-008,
  8.0159e-011, -4.700796e-012, 4.845851e-010, -7.974645e-009,
  -2.475151e-012, -1.377458e-012, 2.437135e-010, 9.211124e-009,
  5.80483e-011, -3.514054e-012, 4.997801e-010, -4.171191e-009,
  -4.789015e-012, -9.645068e-013, 1.761011e-010, 7.839955e-009,
  4.196778e-011, -2.990082e-012, 5.069564e-010, -1.585196e-009,
  -5.260951e-012, -6.037321e-013, 1.138369e-010, 6.52714e-009,
  3.038299e-011, -2.004317e-012, 4.51454e-010, 1.537103e-010,
  -4.860984e-012, -3.502233e-013, 2.678637e-011, 5.298373e-009,
  2.202657e-011, -9.555051e-013, 2.447162e-010, 1.14749e-009,
  -3.956333e-012, -1.444934e-013, -4.67014e-011, 4.20028e-009,
  1.60271e-011, -1.346015e-014, 9.520495e-011, 1.819845e-009,
  -2.945642e-012, -1.033407e-013, -5.606798e-011, 3.255654e-009,
  1.172659e-011, 5.614317e-014, 9.140683e-011, 2.180401e-009,
  -1.993513e-012, -1.420669e-013, -4.086042e-011, 2.44781e-009,
  8.651827e-012, -2.184647e-013, 1.122908e-010, 2.291712e-009,
  -1.152061e-012, -1.105904e-013, -1.984695e-011, 1.834132e-009,
  6.443521e-012, -1.207097e-013, 3.600868e-011, 2.226662e-009,
  -4.030733e-013, -1.640967e-013, 1.189221e-011, 1.364811e-009,
  4.92898e-012, -6.006657e-014, 8.876035e-011, 2.25896e-009,
  1.348168e-013, -2.061452e-014, -7.309407e-011, 8.463812e-010,
  3.874403e-012, -3.240642e-014, 2.109272e-011, 2.033543e-009,
  5.3137e-013, -8.408332e-014, -2.027151e-011, 6.018057e-010,
  3.08698e-012, -7.496643e-014, 1.418742e-012, 1.818797e-009,
  7.889236e-013, -1.109751e-013, -2.087747e-011, 3.534382e-010,
  2.642339e-012, -7.064724e-014, -6.745863e-012, 1.64688e-009,
  9.607634e-013, -2.168681e-014, -9.835631e-013, 2.139183e-010,
  2.267779e-012, 6.166144e-014, 5.995857e-012, 1.465069e-009,
  1.118341e-012, 1.017795e-014, -6.886021e-013, 7.455424e-011,
  2.005356e-012, 5.600199e-015, -2.306482e-011, 1.280499e-009,
  1.187108e-012, -3.197527e-014, -1.403617e-012, -3.718921e-012,
  1.807858e-012, 2.249393e-014, -2.673173e-012, 1.148689e-009,
  1.22496e-012, 3.843323e-014, 1.299065e-011, -4.973894e-011,
  1.652144e-012, -2.050924e-014, -2.361161e-011, 9.67078e-010,
  1.222191e-012, 1.614267e-015, 1.909423e-011, -9.74678e-011,
  1.540309e-012, 2.05924e-014, -1.409442e-011, 8.692258e-010,
  1.17194e-012, -4.981539e-014, -7.464866e-012, -1.395508e-010,
  1.444699e-012, -2.217324e-014, 1.532392e-011, 7.883346e-010,
  1.127552e-012, -2.320003e-015, 2.030727e-011, -1.090925e-010,
  1.36891e-012, 3.539216e-014, 1.281149e-011, 6.75932e-010,
  1.061692e-012, 2.83126e-014, 9.485453e-012, -1.386952e-010,
  1.286977e-012, 3.368452e-014, -1.364666e-011, 5.778004e-010,
  9.869469e-013, -2.233786e-014, 7.0174e-012, -1.344557e-010,
  1.225059e-012, 5.305836e-014, -2.179925e-011, 5.023298e-010,
  9.294074e-013, -1.933389e-014, -7.997498e-012, -1.645722e-010,
  1.148536e-012, 3.108838e-014, -3.308587e-011, 4.254713e-010,
  8.86725e-013, -1.906275e-014, 3.101111e-011, -1.005164e-010,
  1.084379e-012, 2.837677e-014, -8.742868e-012, 4.003808e-010,
  7.892259e-013, -7.533407e-014, -3.147952e-011, -1.742601e-010,
  1.008326e-012, -8.063527e-014, 9.712175e-012, 3.657903e-010,
  7.220138e-013, -8.134751e-014, 5.069939e-012, -7.258139e-011,
  9.412735e-013, -7.801142e-014, 1.87245e-011, 3.115414e-010,
  6.576119e-013, -2.904648e-014, -4.207835e-011, -1.416275e-010,
  8.66874e-013, -1.421839e-014, 3.976364e-011, 3.120056e-010,
  5.928542e-013, 3.022994e-014, 5.351974e-012, -8.674414e-011,
  8.684767e-013, 1.887022e-013, 3.933496e-011, 2.648208e-010,
  6.662239e-013, -2.502371e-014, 1.260173e-011, -8.110269e-011,
  8.961436e-013, -1.097614e-013, 2.502163e-011, 2.552082e-010,
  5.26681e-013, -2.119729e-014, 3.214558e-011, -1.080009e-011,
  7.854245e-013, 8.791902e-014, -1.210211e-011, 2.053196e-010,
  4.50546e-013, -5.438869e-014, 2.640404e-012, -1.939657e-011,
  7.337076e-013, 4.81456e-014, 2.121166e-011, 2.360414e-010,
  4.176633e-013, -1.624801e-014, 1.387832e-011, -6.809724e-012,
  6.656934e-013, 7.211662e-014, 3.108618e-011, 2.180527e-010,
  3.602815e-013, 4.837297e-014, 1.603864e-011, -9.351899e-012,
  5.806896e-013, 2.352725e-014, -1.443846e-011, 1.294815e-010,
  3.709123e-013, 1.562748e-014, 1.652513e-011, -6.297945e-012,
  5.920101e-013, -1.097641e-014, 1.812218e-011, 1.424648e-010,
  3.512671e-013, -1.164464e-014, -2.087708e-012, -2.606884e-011,
  5.446225e-013, -3.184132e-014, 3.713304e-011, 1.766994e-010,
  3.178869e-013, -3.912513e-014, -1.378426e-011, -4.267522e-011,
  5.098719e-013, -5.357664e-014, 2.534984e-011, 1.530782e-010,
  3.630756e-013, -2.39741e-014, -1.640435e-011, -4.404663e-011,
  4.939003e-013, -1.938338e-014, 5.739647e-013, 1.064982e-010,
  3.232627e-013, 6.788679e-015, -9.065791e-012, -3.54177e-011,
  4.674049e-013, -3.726625e-015, -1.4918e-011, 6.824442e-011,
  2.52142e-013, -4.539363e-014, 1.178293e-012, -8.009268e-012,
  4.343954e-013, -4.195054e-014, 1.054097e-011, 9.998687e-011,
  2.675939e-013, -1.348121e-014, 5.169055e-011, 3.646932e-011,
  4.274255e-013, -4.100714e-014, -1.701138e-011, 5.513977e-011,
  2.357269e-013, -1.214218e-014, 4.596953e-011, 5.69286e-011,
  3.80475e-013, -1.612684e-014, 2.187666e-011, 1.096075e-010,
  1.96488e-013, -5.890887e-014, -2.389025e-011, -5.467434e-011,
  3.896293e-013, -1.005813e-014, 1.297661e-011, 1.104909e-010,
  2.276485e-013, 7.763251e-014, 3.296921e-011, 8.225611e-012,
  3.494079e-013, -4.515839e-014, -9.182284e-011, -6.214972e-011,
  2.212229e-013, -1.965321e-015, -2.565794e-011, -7.201576e-011,
  3.100018e-013, -7.341865e-014, -4.481988e-011, 2.648664e-011,
  1.856489e-013, -5.862233e-014, -2.310104e-011, -2.671944e-011,
  2.841682e-013, 5.198523e-014, 4.698023e-011, 1.47535e-010,
  2.773009e-013, -2.804962e-014, 1.255017e-011, 8.45077e-012,
  3.864285e-013, -5.017348e-015, 3.093939e-011, 8.835128e-011,
  1.491383e-013, 2.682901e-014, 2.103924e-011, -6.404e-013,
  2.492859e-013, -8.115915e-014, -5.673392e-013, 4.918721e-011,
  1.634117e-013, -4.640915e-014, 1.14664e-011, 7.178279e-012,
  2.322481e-013, -9.988641e-014, -3.399311e-011, -5.81873e-012,
  1.726467e-013, 6.087517e-014, 3.208926e-011, 3.841426e-011,
  2.447013e-013, -1.010603e-014, -1.631162e-012, 2.927509e-011,
  9.339311e-014, -5.392236e-014, -3.100216e-012, 8.980253e-012,
  1.714315e-013, -4.040185e-014, 3.100184e-011, 8.89353e-011,
  1.422783e-013, -3.641111e-014, 9.707517e-012, 5.094791e-012,
  2.233115e-013, -7.037183e-014, 2.057174e-011, 5.352806e-011,
  1.31653e-013, -6.235993e-014, 1.695804e-012, 1.076918e-011,
  2.122883e-013, -1.063585e-013, 1.31272e-011, 4.131749e-011,
  1.248811e-013, -5.64725e-014, 5.476472e-012, 8.358409e-012,
  2.045706e-013, -4.394152e-015, 2.135261e-011, 7.0976e-011,
  1.807499e-013, -6.989676e-014, -2.703008e-011, -6.463499e-011,
  2.03247e-013, -1.074158e-013, 3.693999e-012, 5.447486e-011,
  1.359374e-013, -1.20902e-014, -1.415621e-011, -3.891047e-011,
  1.817748e-013, -8.45139e-014, 1.997295e-012, 3.69023e-011,
  1.080098e-013, -3.66385e-014, 8.936413e-012, 7.546782e-013,
  1.831307e-013, -6.410196e-014, 8.608886e-012, 3.413969e-011,
  1.028379e-013, -5.548409e-014, 2.721308e-012, -5.812274e-012,
  1.630459e-013, -5.053942e-014, 1.1952e-011, 4.591035e-011,
  1.063368e-013, -1.603337e-014, -5.051311e-013, 1.362302e-012,
  1.684676e-013, -1.170197e-015, 1.583816e-011, 5.761039e-011,
  9.000975e-014, -7.747465e-014, -2.342368e-011, -3.268457e-011,
  1.430519e-013, -8.718567e-014, 1.229692e-011, 5.991537e-011,
  8.879222e-014, -4.173666e-014, 1.733593e-011, 2.957368e-011,
  1.475223e-013, -2.659948e-014, 2.538445e-011, 6.875039e-011,
  1.045882e-013, -3.36879e-014, 1.211058e-012, -1.546415e-011,
  1.369867e-013, -3.839561e-014, 7.807525e-012, 3.340951e-011,
  9.257828e-014, 6.007447e-014, -2.411926e-011, -6.844322e-011,
  1.41388e-013, -7.529508e-014, -1.86167e-011, -1.562491e-011,
  1.262712e-013, -1.783803e-014, -5.464067e-011, -8.359321e-011,
  2.035596e-013, -2.760669e-015, 4.339672e-011, 1.024409e-010,
  8.287803e-014, 2.671923e-015, 1.638306e-011, 2.540134e-011,
  1.275581e-013, 5.971546e-014, -1.834459e-012, 1.418187e-011,
  7.105431e-014, -1.562754e-014, 4.217949e-012, -1.222961e-011,
  1.329437e-013, -6.870108e-014, 5.624829e-012, 4.163779e-011,
  6.746124e-014, -1.014082e-014, 5.229158e-011, 3.901479e-011,
  1.432071e-013, -2.970362e-014, -7.062531e-011, -5.410783e-011,
  2.754443e-014, -8.120922e-014, 7.995377e-011, 9.965694e-011,
  5.668829e-014, -2.326444e-014, -1.922295e-011, 4.186326e-011,
  4.317857e-014, 1.708437e-013, -9.960621e-011, -1.804298e-010,
  1.210923e-013, -2.308718e-014, -7.138713e-011, -7.398199e-011,
  7.715177e-014, -4.299688e-014, -2.887637e-011, -3.149567e-011,
  7.410747e-014, 1.674894e-013, 4.519541e-011, 1.075113e-010,
  1.884286e-013, -1.886214e-013, -7.291253e-011, -8.163015e-011,
  4.224586e-014, 9.300483e-014, -6.9559e-013, 8.019752e-011,
  -3.681847e-014, 2.217473e-014, 6.195513e-011, 6.120066e-011,
  3.372505e-013, -4.137506e-014, 1.167653e-010, 1.676093e-010,
  -1.60518e-013, 2.643795e-014, -2.891243e-011, -5.432201e-011,
  1.051309e-013, -2.925367e-014, 1.673413e-010, 2.096588e-010,
  -1.450923e-013, 2.40619e-014, 4.014289e-011, 4.429124e-011,
  1.099863e-013, -7.427833e-014, 1.015086e-010, 1.206752e-010,
  -1.859652e-013, -7.489866e-015, -6.66131e-011, -7.036539e-011,
  1.966049e-013, 1.034944e-014, 1.270212e-010, 1.766147e-010,
  -9.89294e-014, 5.729251e-014, -2.966884e-012, 2.24357e-011,
  9.435165e-014, 4.902475e-014, 4.656589e-011, 6.350309e-011,
  -1.002514e-013, -4.614431e-014, 6.135665e-012, -7.255112e-012,
  2.350046e-013, -5.334907e-014, 1.806393e-010, 2.308982e-010,
  4.893486e-014, -2.757324e-014, -1.196825e-013, -3.754086e-011,
  -3.435916e-014, 4.073975e-014, 1.00266e-010, 1.816669e-010,
  -1.938026e-014, 4.03016e-014, -3.020987e-011, -1.390631e-011,
  1.073384e-013, 2.56623e-014, 1.482584e-011, 6.618538e-011,
  4.468595e-014, 4.50852e-015, -4.602554e-011, -8.525426e-011,
  1.682964e-014, -5.184179e-014, -4.845026e-011, -5.050305e-011,
  -4.981487e-014, -2.870525e-014, -8.196208e-011, -1.353677e-010,
  2.098866e-013, -2.970338e-014, -6.029864e-012, -1.536259e-012,
  6.372376e-014, -5.222327e-014, 5.619039e-011, 6.30152e-011,
  1.131565e-013, -1.899644e-014, 1.365251e-011, 5.075299e-011,
  4.154464e-014, 1.038427e-014, 1.269566e-011, -3.224331e-013,
  9.972264e-014, -2.200899e-014, 3.500971e-011, 7.21667e-011,
  3.757507e-014, -2.191353e-014, 4.369822e-012, 6.779706e-012,
  1.273163e-013, -6.1378e-014, 6.272712e-011, 9.121441e-011,
  1.867291e-015, 2.232339e-014, 7.534061e-012, 9.299238e-012,
  1.02094e-013, -3.991846e-014, 2.005688e-011, 1.569282e-011,
  5.87658e-015, -7.690325e-014, -2.41987e-011, -5.184779e-011,
  5.157769e-014, -4.672981e-014, 5.469005e-011, 9.303462e-011,
  1.340084e-014, 3.590219e-015, -2.166295e-011, -2.646441e-011,
  2.723548e-014, -1.701246e-014, -1.124132e-011, -1.122094e-011,
  4.316252e-014, -1.801776e-014, -1.792658e-011, -2.747806e-011,
  3.116162e-014, -4.602855e-015, -1.445769e-011, -1.153695e-011,
  3.685312e-014, 2.560008e-015, -2.130082e-011, -2.0985e-011,
  1.966879e-014, 1.808886e-016, -2.256147e-011, -2.577796e-011,
  5.421746e-014, -1.475453e-014, -2.11252e-011, -2.573802e-011,
  2.791584e-014, -1.807316e-014, -8.314785e-012, -3.777436e-012,
  3.1514e-014, -2.830795e-014, -5.551307e-012, -9.998764e-012,
  4.652174e-014, -2.360819e-014, 1.363694e-011, 2.29415e-011,
  2.274889e-014, -3.36788e-014, -4.297677e-014, -2.165712e-011,
  4.801308e-014, -2.562297e-014, 1.138031e-011, 9.723948e-012,
  5.473397e-014, -2.825636e-014, -6.48294e-012, -2.115063e-011,
  -6.151335e-016, -3.435262e-014, 1.35138e-011, 8.028912e-012,
  4.051927e-014, 1.975733e-014, 1.155043e-011, 2.121579e-011,
  1.23473e-014, 1.045709e-015, -9.700734e-012, -1.931919e-012,
  4.953945e-014, 7.752527e-014, -3.257388e-012, -2.942269e-011,
  6.13883e-014, -6.699035e-014, -2.453548e-011, -1.90714e-011,
  3.062145e-014, -2.291384e-014, -1.158449e-011, -3.013443e-011,
  7.847606e-014, -3.042061e-014, -3.188539e-012, 1.467606e-011,
  6.344734e-015, -5.016636e-014, 9.135444e-012, 9.199179e-012,
  9.038018e-014, -2.149971e-014, 3.002908e-011, 5.213037e-011,
  5.712253e-014, 3.55851e-014, 4.873004e-011, 6.135454e-011,
  1.157223e-013, -4.239327e-015, -1.74382e-011, -3.940936e-011,
  5.66908e-014, 3.29453e-014, 9.951852e-012, -5.912218e-012,
  5.043607e-014, -2.913768e-014, -1.555359e-011, -3.812699e-011,
  1.314677e-014, -2.370397e-014, -2.407361e-011, -1.993377e-011,
  -2.0905e-014, -8.22646e-015, 5.492324e-011, 7.838199e-011,
  1.461758e-014, -7.857758e-015, -8.544667e-011, -9.987898e-011,
  -4.577722e-014, 1.794161e-014, 8.632894e-011, 1.225784e-010,
  1.594321e-013, -3.567776e-014, 9.627667e-011, 1.286194e-010,
  -1.166079e-013, -2.479953e-014, 1.623088e-010, 2.408564e-010,
  1.339004e-013, -2.371534e-014, 4.356107e-011, 3.049308e-011,
  3.229867e-013, -6.679771e-014, 4.763917e-011, 1.12296e-010,
  3.662086e-013, -6.442715e-014, 9.531688e-011, 1.466955e-010,
  -1.416237e-014, 1.128728e-014, -4.855317e-011, -3.022298e-011,
  3.248316e-013, -4.854856e-014, 1.690628e-010, 2.046215e-010,
  1.462821e-013, -4.947569e-014, 3.508428e-011, 7.204906e-011,
  5.827516e-014, -2.971978e-014, 1.32799e-010, 1.627558e-010,
  2.039288e-013, -5.262626e-014, 6.023905e-012, 4.883049e-012,
  -1.599514e-013, 1.578011e-014, -7.397663e-011, -1.01464e-010,
  -1.130902e-014, -3.193895e-014, 8.352821e-011, 9.802302e-011,
  -3.704166e-013, 1.445682e-013, 7.846202e-012, -3.521351e-011,
  1.736239e-013, -1.115809e-013, 1.989057e-010, 2.222449e-010,
  -1.114082e-013, -5.507506e-014, -6.360835e-011, -1.146517e-010,
  1.048869e-013, -8.755437e-014, -3.961663e-011, -6.32355e-011,
  -3.333033e-014, -1.059581e-013, 1.155523e-010, 1.073216e-010,
  3.848828e-014, -2.164492e-016, 1.282227e-010, 1.820512e-010,
  1.390653e-013, -1.408366e-014, 1.112031e-010, 1.402123e-010,
  -1.036588e-013, 4.891749e-014, 5.829615e-011, 8.695384e-011,
  3.130848e-014, -1.672378e-014, -1.190708e-010, -1.11319e-010,
  -3.942981e-013, 1.614044e-013, -1.246783e-010, -1.534585e-010,
  8.396071e-014, -3.696544e-014, 9.964272e-011, 1.492843e-010,
  -1.027945e-013, 1.690921e-014, -1.979685e-011, -2.317605e-011,
  -5.114113e-014, -7.899538e-014, 3.205983e-012, 5.400504e-011,
  -1.554255e-013, 9.20987e-014, 4.439046e-011, 6.726775e-011,
  -1.715644e-014, -6.545486e-014, 4.678561e-011, 4.35806e-011,
  -7.578948e-015, -1.023169e-013, 3.154477e-011, -8.951317e-012,
  -3.9125e-014, -4.62102e-014, 1.100818e-012, 1.53658e-012,
  1.06379e-013, -8.271987e-014, 5.475056e-011, 3.518804e-011,
  -5.83156e-014, -4.27906e-014, 1.237861e-011, 1.503376e-011,
  1.013762e-013, -3.920645e-014, 5.300696e-011, 6.730257e-011,
  1.547503e-013, -4.424942e-014, -8.071777e-012, -1.59836e-011,
  6.70204e-014, -2.964891e-014, 2.735105e-011, 5.868354e-011,
  9.619833e-014, -4.623631e-014, -7.785383e-012, -1.142747e-011,
  -9.295738e-015, -1.49907e-014, -3.299589e-012, 5.467535e-012,
  9.521649e-014, -2.005158e-014, 9.0306e-012, 3.640658e-011,
  -6.692676e-014, 2.36522e-014, -5.586099e-011, -6.794197e-011,
  -1.349661e-014, 8.249538e-015, -3.701095e-011, -4.744299e-011,
  4.386062e-014, -1.40033e-014, -4.587056e-012, -9.027903e-012,
  -4.34825e-014, 1.463116e-014, -6.527858e-011, -7.46558e-011,
  4.791797e-015, -8.275532e-015, 2.7169e-011, 2.173017e-011,
  -9.803819e-014, -2.856435e-014, -2.991756e-011, -5.372488e-011,
  4.590219e-014, -3.274025e-014, 3.977473e-011, 4.413418e-011,
  -5.597377e-015, 1.705896e-014, 1.293459e-011, 3.754243e-011,
  9.382557e-015, 4.966006e-014, 2.891051e-011, 3.519965e-011,
  -1.105643e-013, -1.908061e-014, 4.465269e-012, 2.277701e-011,
  9.272758e-014, 5.243261e-014, 5.314967e-011, 6.921466e-011,
  -1.270578e-013, 5.932197e-014, -3.589831e-011, -5.7504e-011,
  1.3963e-013, -1.059856e-013, 2.597997e-011, -1.078084e-012,
  -3.444364e-014, 4.381831e-014, -7.365442e-013, -3.505735e-012,
  -3.093182e-014, 2.75868e-014, 2.290466e-011, 1.969329e-011,
  1.017197e-013, -5.431601e-014, -5.631916e-012, 1.119859e-011,
  3.109028e-014, -4.187038e-014, -7.735466e-011, -1.135911e-010,
  2.392987e-013, 4.650902e-015, 9.080239e-012, 4.341326e-011,
  2.114778e-014, 2.261171e-014, -9.662819e-012, -1.648645e-011,
  2.571016e-014, -1.577371e-014, -3.747434e-011, -5.789404e-011,
  1.509187e-013, 3.395146e-014, 2.868669e-011, 4.97986e-011,
  -5.959939e-014, 6.017338e-014, -1.024875e-010, -1.178492e-010,
  -2.900258e-013, 1.012446e-013, -9.604011e-011, -1.522253e-010,
  -2.282091e-013, -1.359976e-014, -1.255133e-010, -1.328991e-010,
  -1.719092e-013, 2.116283e-014, 5.386152e-013, -6.740132e-012,
  -2.60707e-013, 9.353988e-014, -5.174547e-011, -1.019236e-010,
  7.104828e-014, -3.531687e-014, 1.247749e-010, 1.367992e-010,
  -1.061503e-013, 5.617428e-014, -1.167754e-010, -1.470507e-010,
  3.300101e-015, 6.00904e-015, 6.524065e-011, 7.864433e-011,
  1.56342e-013, -5.050383e-014, 4.840089e-011, 6.768191e-011,
  8.714419e-014, -2.03163e-014, 4.251158e-011, 8.554515e-011,
  1.220721e-013, 5.997668e-014, -3.310023e-011, -2.634559e-011,
  -2.614418e-014, 6.568612e-014, -4.784281e-011, -6.497897e-011,
  -6.224613e-014, 3.161015e-014, -3.24542e-011, -3.596437e-011,
  2.244908e-014, -6.923587e-015, -3.204507e-011, -7.990897e-011,
  -6.192552e-015, -2.088284e-014, -3.427351e-011, -2.730939e-011,
  -1.039095e-013, -3.332088e-015, -3.679353e-011, -4.23373e-011,
  8.879751e-014, -3.644307e-014, -1.247337e-011, 1.309962e-011,
  -1.343958e-013, 6.888727e-014, -1.357941e-011, -1.569093e-011,
  -1.570449e-013, 6.274252e-015, -4.640322e-011, -5.164199e-011,
  -1.782154e-014, 2.659967e-014, -1.559655e-011, -2.278764e-011,
  3.044999e-014, -1.064015e-015, -1.477538e-011, -1.842551e-011,
  5.668711e-014, -1.311133e-014, -2.435145e-011, -6.380569e-012,
  4.255105e-015, -1.77024e-015, -1.787161e-011, -1.693184e-011,
  -7.365934e-015, 6.397028e-014, 1.512124e-011, 3.250478e-011,
  7.353034e-014, -6.108794e-017, -4.283125e-011, -7.594044e-011,
  1.523803e-013, 1.341301e-014, 5.394e-011, 8.653553e-011,
  -6.060332e-014, 6.957009e-015, 3.717717e-011, 5.337254e-011,
  -6.552631e-014, 1.45066e-014, 1.846808e-011, 4.553981e-011,
  5.728367e-015, 5.027274e-014, -2.422696e-011, -2.749085e-011,
  9.382457e-014, -4.992741e-014, -2.411938e-011, -2.518657e-011,
  7.911699e-014, -6.04743e-014, -2.76749e-011, -4.851644e-011,
  4.18036e-014, -9.055315e-014, 9.684946e-012, 2.93697e-011,
  -2.376081e-013, 5.900426e-015, -9.722859e-011, -7.580813e-011,
  -2.438297e-013, 6.013655e-014, 5.475133e-011, 5.844179e-011,
  -2.300432e-013, 2.61841e-014, -6.560707e-011, -8.796753e-011,
  -1.305144e-013, 3.229443e-014, 1.371799e-010, 1.603075e-010,
  -1.399003e-013, 2.187458e-015, -6.725384e-011, -4.215826e-011,
  -7.331858e-014, 7.373413e-014, 1.855729e-011, 1.853082e-011,
  -5.011587e-014, 2.771283e-014, 1.868388e-011, 1.168753e-011,
  5.207138e-014, -5.22245e-014, -5.178597e-011, -8.578962e-011,
  -2.584631e-013, 1.337618e-013, -7.313652e-011, -7.752125e-011,
  -3.378542e-013, 5.394524e-014, -2.215173e-010, -3.510646e-010,
  -2.790685e-013, 1.371981e-014, -1.420624e-010, -1.674025e-010,
  -6.518396e-014, 1.070579e-016, -6.524568e-011, -1.282785e-010,
  -2.507732e-014, 3.986173e-014, 3.81856e-011, 6.771797e-011,
  2.09549e-013, -5.530788e-014, -2.259384e-011, -2.99726e-011,
  -2.619708e-013, 1.098406e-013, -2.155736e-010, -2.253157e-010,
  -2.34139e-013, 6.979085e-014, -1.11682e-010, -1.950032e-010,
  -1.679224e-013, -5.967729e-015, -1.036864e-010, -1.789117e-010,
  2.937298e-014, -1.067905e-013, 5.658955e-011, 7.00839e-011,
  -7.31564e-014, -3.597091e-014, -3.010671e-011, -4.654459e-011,
  -4.891065e-014, 3.007318e-014, 1.236497e-010, 2.195325e-010,
  7.186057e-014, -2.770283e-014, 2.642986e-011, 3.154906e-012,
  6.777427e-015, -4.196401e-014, 1.255864e-010, 1.876021e-010,
  7.927264e-014, 3.985917e-014, 7.798132e-011, 8.70384e-011,
  1.296631e-013, -5.778217e-015, 2.607941e-014, -2.633192e-012,
  -1.164156e-014, 3.16816e-014, 4.956663e-011, 7.311965e-011,
  1.291339e-013, 1.453714e-015, 1.649882e-011, -3.752252e-012,
  5.2355e-014, -2.010771e-015, 8.802584e-011, 1.20338e-010,
  1.565742e-013, -9.980584e-014, 5.195572e-011, 8.609294e-011,
  -5.417854e-014, 7.236992e-014, 4.750268e-011, 5.177717e-011,
  3.508493e-014, -7.673602e-014, -6.096043e-012, -2.811612e-011,
  -1.942114e-013, 7.096215e-014, -2.752776e-011, -4.415927e-011,
  -4.023642e-014, -3.029341e-014, 3.547228e-011, 1.370806e-011,
  1.85392e-014, -1.231473e-013, -5.702549e-011, -9.011757e-011,
  -7.076583e-014, -4.896724e-014, -1.401803e-011, 5.471409e-012,
  2.222701e-014, 2.757793e-014, 3.935378e-011, 4.065319e-011,
  -3.146244e-014, -7.688813e-014, -9.349234e-012, -2.433673e-011,
  -1.562779e-013, 1.400852e-013, -1.671088e-011, -9.764828e-012,
  -7.987679e-014, 1.398968e-014, 2.809338e-011, -1.227695e-011,
  -4.053154e-014, 3.249677e-014, -8.148713e-011, -9.589166e-011,
  -1.183569e-013, 3.358315e-014, 4.937252e-011, 4.325341e-011,
  -2.591432e-015, 9.980782e-014, -6.578643e-011, -1.118131e-010,
  -5.602063e-014, -1.539306e-014, 9.013282e-012, -1.467515e-011,
  3.335511e-013, -1.784009e-014, -4.937729e-012, -1.518875e-011,
  -1.117477e-013, 3.163492e-014, -1.626168e-011, 9.131112e-012,
  4.381137e-013, -1.350612e-013, -6.131735e-011, -1.217634e-010,
  -5.409959e-014, -1.877131e-014, -2.007212e-012, 3.417972e-011,
  2.184815e-013, 1.743814e-014, 8.570133e-011, 9.779417e-011,
  -4.12719e-014, 5.50462e-014, -9.626474e-011, -1.438256e-010,
  -3.539476e-014, -2.717876e-014, 5.272441e-011, 1.719037e-011,
  1.752013e-013, -9.740172e-014, 1.24191e-010, 1.818289e-010,
  7.72768e-014, 1.610188e-014, -2.147379e-012, -4.297312e-011,
  -1.77892e-014, -5.79639e-014, 8.07877e-011, 1.161125e-010,
  -1.267207e-013, 7.237357e-014, -1.121899e-011, -1.747965e-012,
  -2.447863e-013, -9.866008e-016, -7.069985e-011, -3.932563e-011,
  -1.277026e-013, 3.031049e-014, -1.80977e-011, 3.057679e-011,
  -6.187482e-014, 3.091609e-014, -1.337047e-010, -1.782685e-010,
  -9.408992e-014, -3.713919e-014, 1.011696e-010, 1.585123e-010,
  2.426064e-013, 1.385741e-014, 2.603901e-010, 3.555952e-010,
  -5.948461e-014, -1.359892e-014, -5.754704e-011, -1.440834e-010,
  -6.375788e-014, -1.672173e-013, 1.486391e-010, 1.810117e-010,
  -3.213728e-013, 2.629992e-014, 6.478799e-011, 5.559055e-011,
  1.365793e-013, 6.127987e-014, 2.264965e-010, 3.299744e-010,
  1.378294e-014, -2.837222e-015, 1.261524e-012, -1.035538e-012,
  2.078838e-014, 4.029087e-015, -6.397146e-012, 1.656592e-012,
  1.567319e-014, -2.388348e-015, -3.080767e-011, -1.690827e-011,
  -1.179007e-014, 6.498934e-015, -3.654506e-011, -2.105845e-011,
  -6.58631e-015, 3.135034e-015, 1.680419e-012, 1.948218e-012,
  -9.723474e-014, 1.845269e-014, -7.860077e-012, -7.03075e-014,
  1.415725e-014, 1.119323e-014, 6.624948e-012, 4.661597e-012,
  3.140948e-015, 2.973391e-015, -1.700113e-011, -5.820901e-012,
  1.332695e-014, 9.336707e-016, 2.991008e-012, 3.979599e-012,
  2.527287e-014, 3.34532e-015, -1.894028e-012, 8.429214e-012,
  2.254805e-014, 1.484643e-015, -2.869967e-012, 1.009843e-011,
  1.677667e-014, 5.820186e-015, 1.546436e-011, 1.360812e-011,
  9.96661e-014, -6.017975e-015, 1.391811e-011, 1.29643e-011,
  1.90361e-014, 7.765893e-015, -1.06817e-011, -3.022266e-012,
  1.655728e-014, 4.160597e-015, 1.510515e-011, 1.702724e-011,
  2.207368e-014, 1.392302e-014, 2.382904e-013, 8.443337e-012,
  1.544681e-014, 2.233157e-015, -1.523056e-011, -3.245293e-012,
  2.105726e-014, 1.601591e-015, -1.593966e-011, 6.530868e-014,
  8.9753e-015, -3.94114e-014, -1.942865e-011, -6.237187e-012,
  1.640116e-014, -5.502081e-014, -1.308151e-011, 4.900884e-013,
  -4.632738e-014, 1.514751e-014, -8.917409e-013, -8.94232e-013,
  -2.105966e-014, 1.946926e-014, -1.935452e-012, 1.01787e-011,
  4.479831e-015, 3.848445e-015, -1.82875e-012, -2.779155e-012,
  2.429367e-014, 1.561689e-015, -1.227877e-012, 6.674179e-012,
  1.501807e-014, 1.03905e-015, 5.220523e-012, -6.185482e-013,
  2.921914e-014, 8.398494e-015, 4.629714e-013, 9.09189e-012,
  1.541919e-014, 4.906612e-015, 4.590084e-012, -9.03977e-013,
  2.578399e-014, 3.440668e-015, 1.744218e-013, 9.739386e-012,
  2.239279e-014, -1.095813e-015, -4.81798e-012, -5.396062e-012,
  2.825621e-014, 2.730833e-015, 2.641571e-013, 8.67123e-012,
  2.171261e-014, 1.855003e-015, -4.138021e-012, -7.518273e-012,
  2.418338e-014, 2.202274e-015, 4.745442e-012, 1.317618e-011,
  1.800189e-014, 1.598378e-015, -5.45337e-012, -5.14356e-012,
  2.636173e-014, -8.110571e-018, -3.701383e-012, 2.185363e-012,
  2.529451e-014, 1.648261e-015, -6.158781e-013, -7.486187e-013,
  3.61019e-014, -5.062797e-016, 5.540287e-013, 1.13782e-011,
  2.013036e-014, -1.204817e-014, 4.25596e-013, -4.6716e-013,
  3.283529e-014, -4.917006e-015, 2.153742e-013, 9.530252e-012,
  1.83515e-014, -5.860154e-015, 1.41633e-012, 8.055251e-014,
  3.255026e-014, -3.086488e-015, -9.469464e-012, -3.884088e-012,
  2.479045e-014, 1.866266e-015, -7.234001e-013, -1.69648e-012,
  3.436011e-014, 4.243333e-015, -7.290127e-012, 2.609305e-012,
  2.205907e-014, 5.080888e-015, -7.141239e-012, -3.132389e-012,
  3.699443e-014, 3.893627e-016, -2.651515e-012, 1.135765e-011,
  3.372178e-014, -1.295929e-015, 1.767503e-012, 9.195876e-013,
  3.805405e-014, 1.720419e-016, 2.365629e-012, 1.079814e-011,
  1.027992e-013, -1.1706e-014, -5.915258e-012, -8.325297e-012,
  4.589558e-014, -2.510504e-015, 1.582846e-012, 5.350278e-012,
  2.364375e-014, 2.524167e-015, -3.213366e-012, -1.511084e-012,
  3.235478e-014, -6.790105e-015, -6.34607e-013, 1.170416e-011,
  2.719693e-014, -9.816494e-016, -5.223359e-012, -5.187019e-012,
  4.095033e-014, -4.735122e-015, -1.402712e-011, -1.314014e-012,
  2.570378e-014, 4.050051e-015, -7.57947e-013, -2.224134e-012,
  4.058704e-014, -1.031855e-014, -6.129016e-012, 5.877326e-012,
  -4.153333e-014, 1.413448e-014, 4.915701e-012, -1.348161e-012,
  -3.812008e-014, 1.586022e-015, 1.18081e-011, 2.305577e-011,
  1.726892e-014, -7.755132e-016, 1.470992e-013, 1.262422e-012,
  3.53621e-014, -1.269162e-014, -6.3355e-015, 1.380847e-011,
  2.524923e-014, 5.759102e-016, -2.18925e-012, 3.769276e-013,
  4.387952e-014, -5.898973e-015, -6.644654e-012, 5.327583e-012,
  2.687546e-014, -5.371779e-015, 1.737802e-012, -1.87951e-012,
  4.633169e-014, -4.634839e-015, 5.730524e-012, 1.187632e-011,
  3.656251e-014, -5.855381e-016, -8.230887e-012, -1.148143e-011,
  4.798274e-014, -6.085197e-015, 5.770525e-012, 1.210448e-011,
  3.317569e-014, -6.061668e-015, -6.432768e-012, -1.028331e-011,
  4.21173e-014, -2.253601e-015, 8.516881e-012, 1.627187e-011,
  2.134677e-014, -1.710432e-015, 2.81891e-012, 5.033776e-012,
  4.10222e-014, 8.343697e-016, -1.752274e-013, 6.38425e-012,
  3.01744e-014, -2.321868e-015, 6.835141e-012, 3.416714e-012,
  5.314873e-014, 3.445905e-016, -7.775619e-013, 1.36505e-011,
  1.034568e-013, -1.467981e-014, -2.886371e-012, -5.10801e-012,
  4.933436e-014, -5.153968e-015, -9.249592e-012, 5.068492e-012,
  1.229554e-013, -1.599127e-014, 1.375945e-011, 1.532111e-011,
  4.088892e-014, -3.517176e-015, -5.554531e-013, 1.384947e-011,
  4.115418e-014, -7.170133e-015, -4.787641e-012, -7.844188e-012,
  5.642009e-014, -6.445053e-015, 3.019379e-012, 1.80187e-011,
  3.764552e-014, -5.337406e-015, -1.0571e-012, -3.91034e-012,
  5.601348e-014, -3.187358e-015, 6.820102e-013, 1.655315e-011,
  3.451847e-014, -4.253901e-015, 3.360669e-013, -4.270102e-012,
  4.921152e-014, 1.497868e-016, 1.677186e-013, 1.862411e-011,
  -5.705317e-015, 4.944659e-015, 1.449248e-012, -3.478044e-012,
  2.590172e-014, 6.737239e-015, -3.365987e-013, 1.824343e-011,
  3.542992e-014, 3.686637e-016, 9.626739e-012, 6.188081e-012,
  7.177072e-014, -6.946709e-016, -1.559004e-012, 1.50407e-011,
  3.919621e-014, 3.555044e-015, 2.909228e-012, 3.27772e-012,
  6.681649e-014, 1.931295e-015, 5.275093e-012, 1.779467e-011,
  4.37848e-014, 3.072908e-015, 1.225488e-012, -2.23116e-012,
  7.053655e-014, 4.084043e-015, 5.141063e-012, 2.219808e-011,
  5.129344e-014, 2.176235e-015, -8.802952e-013, -4.34435e-012,
  1.70107e-013, -1.130354e-014, -3.595009e-012, 1.758204e-011,
  5.783655e-014, 2.437517e-016, 3.943284e-012, -1.348116e-012,
  7.771378e-014, 9.767349e-015, 4.020506e-012, 2.300941e-011,
  4.309914e-014, 1.662243e-014, 6.587048e-012, 6.57503e-012,
  7.96587e-014, 2.597947e-014, -1.135634e-012, 1.744022e-011,
  4.693576e-014, 1.524778e-014, -2.450565e-012, -5.607298e-012,
  7.873401e-014, 1.599062e-014, 9.510484e-013, 2.210133e-011,
  1.405493e-014, 2.204917e-014, -9.793103e-013, -4.603015e-012,
  1.920252e-013, -5.070018e-014, -2.025243e-012, 1.882538e-011,
  5.07342e-014, 8.914751e-015, -1.83312e-012, -8.121992e-012,
  9.849466e-014, 1.387518e-014, 1.447479e-011, 3.668418e-011,
  5.934082e-014, 1.19755e-014, 4.690768e-012, -9.344318e-013,
  8.613732e-014, 1.306823e-014, -7.104143e-012, 2.227099e-011,
  6.273323e-014, 1.155789e-014, -3.305039e-013, -5.521414e-012,
  8.855971e-014, 1.434839e-014, -5.868877e-012, 2.348206e-011,
  1.504518e-014, 1.042415e-014, -1.243749e-012, -3.091132e-012,
  7.371296e-014, 1.692415e-014, 2.68865e-013, 2.797269e-011,
  2.560177e-014, 1.073914e-014, 6.455343e-012, 3.617791e-012,
  9.04532e-014, 9.884202e-015, -2.700289e-012, 2.729338e-011,
  6.808973e-014, 6.591033e-015, 3.962743e-014, -6.080126e-012,
  1.061542e-013, 1.080418e-014, -2.69972e-012, 3.049645e-011,
  7.334978e-014, 6.117859e-015, 1.499151e-012, -6.977701e-012,
  1.097721e-013, 7.085243e-015, 5.426114e-013, 2.971568e-011,
  8.27667e-014, -1.605058e-016, -6.239862e-013, -8.033674e-012,
  1.321699e-013, -3.883454e-015, 2.274292e-013, 2.856582e-011,
  1.139723e-013, 3.860093e-016, -3.435004e-012, -1.022773e-011,
  1.671054e-013, -1.079934e-014, -4.671374e-013, 2.926066e-011,
  8.543348e-014, 7.5779e-015, 1.612627e-012, -5.288533e-012,
  1.210356e-013, -5.879226e-015, 1.097023e-012, 3.429219e-011,
  8.807553e-014, 8.942309e-016, -3.315461e-012, -7.646334e-012,
  1.26676e-013, -4.292044e-015, -2.056812e-013, 3.541294e-011,
  8.924056e-014, -2.519366e-015, 2.375327e-012, -4.595444e-012,
  1.36212e-013, -5.107808e-015, 3.779792e-012, 3.896299e-011,
  8.864478e-014, -2.066988e-015, 1.045876e-012, -6.048593e-012,
  1.404127e-013, -8.332639e-015, 2.105154e-012, 3.894516e-011,
  9.012077e-014, -3.387806e-015, 1.286192e-012, -6.168632e-012,
  1.462366e-013, -6.5813e-015, 1.697274e-012, 3.991518e-011,
  9.736024e-014, -5.408966e-015, 1.251232e-012, -6.658075e-012,
  1.521847e-013, -6.033727e-015, 4.373892e-013, 3.995353e-011,
  9.795193e-014, -5.323009e-015, 7.058813e-013, -8.798074e-012,
  1.598268e-013, -9.023441e-015, -5.509384e-013, 3.924656e-011,
  2.21578e-013, -2.267623e-014, -2.534521e-012, -1.134067e-011,
  1.028484e-013, -3.462857e-015, 9.999251e-014, 3.95005e-011,
  1.172442e-013, -5.592767e-015, 1.307683e-012, -1.042767e-011,
  1.755827e-013, -9.329693e-015, 2.138448e-012, 4.762397e-011,
  1.069278e-013, -2.966646e-014, -1.065405e-012, -1.40168e-011,
  1.857919e-013, -7.61017e-015, 2.13032e-011, 7.78382e-011,
  1.14188e-013, -2.459531e-014, 4.880317e-013, -5.355575e-012,
  1.929327e-013, -4.21435e-015, 1.507025e-011, 7.433684e-011,
  8.184724e-014, 5.492121e-015, -4.049835e-012, -1.649783e-011,
  1.687328e-013, -3.108835e-015, -2.502074e-012, 5.111032e-011,
  1.218307e-013, -3.462939e-015, -3.472715e-012, -1.482936e-011,
  2.056744e-013, -8.3972e-015, 3.037994e-013, 5.712559e-011,
  1.487591e-013, -3.796768e-015, -4.606902e-012, -1.473812e-011,
  2.331136e-013, -7.549222e-015, 1.386738e-011, 7.438044e-011,
  1.492014e-013, -9.145239e-015, 4.408157e-012, -8.152383e-012,
  2.47698e-013, -6.181587e-015, -1.236834e-012, 6.415244e-011,
  1.701555e-013, -8.157496e-015, -6.764118e-013, -1.468213e-011,
  2.160249e-013, -6.573786e-015, 2.499635e-012, 6.996134e-011,
  1.686458e-013, -1.797084e-015, 7.737937e-013, -1.519542e-011,
  2.053e-013, -4.04224e-017, 4.497209e-012, 7.382215e-011,
  1.798036e-013, -1.729885e-015, 2.881181e-013, -1.662846e-011,
  2.745034e-013, -3.158474e-015, 2.826964e-012, 7.707648e-011,
  1.942356e-013, -5.817145e-016, 1.131121e-012, -1.410725e-011,
  2.855514e-013, -3.125892e-015, 1.031456e-012, 8.129746e-011,
  2.027846e-013, -4.260945e-015, 5.86903e-012, -5.985489e-012,
  3.064164e-013, -7.631787e-015, 4.211259e-012, 8.961991e-011,
  2.091389e-013, -9.112535e-015, 6.974222e-012, -5.322924e-012,
  3.317829e-013, -8.637031e-015, 8.064529e-012, 9.450578e-011,
  2.090178e-013, -1.234988e-014, -1.889793e-012, -1.438388e-011,
  3.465168e-013, -7.96426e-015, 1.504817e-011, 1.041209e-010,
  2.285396e-013, -7.50549e-015, 3.438057e-012, -1.785168e-011,
  3.729595e-013, -9.001934e-015, 3.304589e-012, 1.052643e-010,
  2.300195e-013, -3.15411e-015, 4.108656e-012, -2.394653e-011,
  3.935743e-013, -7.793537e-015, 5.929248e-012, 1.170852e-010,
  1.26069e-013, 8.515856e-015, 5.783946e-012, -1.616529e-011,
  3.864339e-013, 7.030683e-015, -6.163585e-012, 1.062082e-010,
  2.834906e-013, 2.960589e-014, 1.056176e-011, -7.987729e-013,
  4.509348e-013, 2.264001e-014, -9.076006e-012, 1.07379e-010,
  2.999464e-013, -9.236848e-015, -2.99054e-012, -2.004439e-011,
  4.775323e-013, -1.512237e-014, -8.311898e-012, 1.210065e-010,
  3.154706e-013, -1.674471e-014, -1.533619e-011, -4.737742e-011,
  5.173122e-013, -3.164085e-014, -5.177462e-012, 1.34159e-010,
  3.545989e-013, -1.733422e-014, 3.52576e-012, -2.377906e-011,
  6.337179e-013, -3.029438e-014, 7.79102e-012, 1.504561e-010,
  3.758256e-013, -1.066249e-014, 4.303325e-012, -2.334297e-011,
  6.118948e-013, -1.793107e-014, 1.262312e-011, 1.649652e-010,
  4.016603e-013, -1.515833e-014, -3.813071e-012, -3.617947e-011,
  6.487861e-013, -2.501275e-014, 9.216005e-012, 1.702607e-010,
  4.373104e-013, -1.538849e-014, -7.314336e-012, -5.398877e-011,
  7.001994e-013, -3.303233e-014, 1.51433e-011, 1.972633e-010,
  4.957178e-013, -5.086299e-014, -5.689844e-012, -4.787164e-011,
  7.10913e-013, -3.599492e-014, 2.004807e-011, 2.017109e-010,
  5.308732e-013, -3.671736e-014, -1.022614e-012, -4.574087e-011,
  7.831879e-013, -3.349994e-014, 2.258183e-011, 2.134701e-010,
  5.665904e-013, -2.263017e-014, 4.948677e-013, -7.167334e-011,
  8.77958e-013, -3.532537e-014, 1.612534e-011, 2.382696e-010,
  6.478677e-013, -1.519884e-014, -1.329983e-011, -8.790497e-011,
  9.499185e-013, -2.32631e-014, 1.552406e-011, 2.485331e-010,
  7.173298e-013, -3.1665e-014, 1.01522e-011, -6.343227e-011,
  1.015091e-012, -1.428689e-014, 1.276327e-011, 2.644701e-010,
  7.717722e-013, -1.641041e-014, 8.466779e-012, -8.500171e-011,
  1.112644e-012, -3.724286e-014, 7.578713e-012, 2.851193e-010,
  8.469572e-013, -2.374259e-014, -1.204607e-012, -1.109593e-010,
  1.192949e-012, -3.836642e-014, 1.203088e-011, 3.251177e-010,
  9.325091e-013, -1.843695e-014, -6.898046e-013, -1.315348e-010,
  1.279284e-012, -2.295259e-014, 7.445145e-012, 3.715842e-010,
  1.030198e-012, -1.655681e-014, -9.643572e-012, -1.575284e-010,
  1.371778e-012, -1.839798e-014, 6.217353e-012, 4.187428e-010,
  1.133291e-012, -1.922821e-014, -2.589674e-012, -1.736904e-010,
  1.468597e-012, -2.237461e-014, 5.140512e-012, 4.794607e-010,
  1.243752e-012, -1.227374e-014, -1.853724e-012, -1.909366e-010,
  1.563319e-012, 1.52947e-016, -1.10163e-012, 5.543849e-010,
  1.356861e-012, -2.577095e-014, 1.284616e-012, -2.017554e-010,
  1.661261e-012, 3.382188e-014, -2.969299e-012, 6.523925e-010,
  1.522078e-012, 1.038124e-014, -6.707945e-012, -2.314748e-010,
  1.782591e-012, 2.74245e-014, -4.554573e-011, 7.095503e-010,
  1.524764e-012, 6.845099e-015, -1.38025e-010, -3.333856e-010,
  1.838859e-012, 1.403202e-014, 6.713775e-011, 9.471582e-010,
  1.585999e-012, 2.063345e-015, 1.893718e-011, -1.727551e-010,
  2.006768e-012, 2.210262e-014, 4.258124e-011, 1.081004e-009,
  1.567799e-012, 1.986989e-014, 3.39061e-011, -1.465519e-010,
  2.188382e-012, 3.434998e-014, 3.327782e-011, 1.256963e-009,
  1.571945e-012, -1.024947e-014, 6.485779e-012, -5.124158e-011,
  2.390894e-012, 9.326919e-015, 7.804538e-012, 1.464233e-009,
  1.457559e-012, -2.303735e-014, 1.449871e-011, 9.388341e-011,
  2.69003e-012, -3.032447e-014, 2.195543e-011, 1.70453e-009,
  1.179053e-012, -4.960852e-014, -2.979136e-011, 2.507079e-010,
  3.098048e-012, -9.966867e-014, 8.296536e-011, 2.027869e-009,
  8.12112e-013, -4.442357e-014, 3.141136e-012, 5.676344e-010,
  3.750635e-012, -9.502889e-014, 5.479725e-011, 2.256337e-009,
  2.475626e-013, -2.246171e-014, 6.551663e-012, 9.746313e-010,
  4.710459e-012, -1.241625e-013, 6.028768e-011, 2.53773e-009,
  -5.01845e-013, -9.638855e-015, 2.518855e-011, 1.527784e-009,
  6.132465e-012, -2.145656e-013, 7.76217e-011, 2.785264e-009,
  -1.511921e-012, -1.24793e-014, 3.500198e-011, 2.25096e-009,
  8.266512e-012, -3.975335e-013, 1.162709e-010, 2.952523e-009,
  -2.741001e-012, -1.233906e-014, 5.704036e-011, 3.174875e-009,
  1.142111e-011, -6.43775e-013, 1.523213e-010, 2.981871e-009,
  -4.195656e-012, -2.962684e-014, 7.877671e-011, 4.308229e-009,
  1.611299e-011, -1.027726e-012, 1.989839e-010, 2.783006e-009,
  -5.707152e-012, -9.95794e-014, 1.151711e-010, 5.740206e-009,
  2.298225e-011, -1.49313e-012, 2.189269e-010, 2.182013e-009,
  -6.898873e-012, -3.124916e-013, 2.075432e-010, 7.432897e-009,
  3.298035e-011, -2.538422e-012, 2.832312e-010, 1.020703e-009,
  -7.045419e-012, -7.727318e-013, 3.05928e-010, 9.290459e-009,
  4.743672e-011, -3.985679e-012, 3.451188e-010, -9.834462e-010,
  -3.811666e-012, -1.496751e-012, 3.486926e-010, 1.125098e-008,
  6.804458e-011, -5.123054e-012, 2.895577e-010, -4.232566e-009,
  3.332196e-012, -3.032945e-012, 3.951622e-010, 1.298188e-008,
  9.879794e-011, -7.000614e-012, 2.398073e-010, -9.348829e-009,
  1.950652e-011, -5.99853e-012, 4.622835e-010, 1.38835e-008,
  1.434278e-010, -1.043397e-011, 2.511992e-010, -1.725744e-008,
  5.268481e-011, -9.945334e-012, 4.525701e-010, 1.281535e-008,
  2.087804e-010, -1.332167e-011, 2.067568e-010, -2.9257e-008,
  1.191369e-010, -1.579603e-011, 3.490539e-010, 7.568632e-009,
  3.04434e-010, -1.590564e-011, 1.764283e-010, -4.700418e-008,
  2.509462e-010, -2.401028e-011, 2.031134e-010, -6.443078e-009,
  4.482029e-010, -1.759105e-011, 2.815023e-010, -7.39132e-008,
  5.130664e-010, -3.594011e-011, 2.091324e-010, -3.834502e-008,
  6.666085e-010, -1.68768e-011, 8.661763e-010, -1.14395e-007,
  1.053035e-009, -6.680951e-011, 1.383861e-009, -1.111804e-007,
  9.984442e-010, -1.608822e-011, 3.26448e-009, -1.773526e-007,
  2.10398e-009, -1.360897e-010, 6.631546e-009, -2.846051e-007,
  1.48289e-009, -1.30317e-011, 8.438824e-009, -2.786517e-007,
  3.090401e-009, -3.158876e-010, 2.671803e-008, -7.415009e-007,
  1.955107e-009, -3.911037e-012, 1.93752e-008, -4.492823e-007,
  -2.228166e-009, -6.43618e-010, 8.918666e-008, -1.875376e-006,
  1.678689e-009, 1.046586e-011, 3.84567e-008, -7.169309e-007,
  -1.218906e-008, -6.794244e-010, 1.482811e-007, -3.236179e-006,
  1.568471e-009, 3.964168e-011, 4.753247e-008, -9.369419e-007,
  -1.423926e-008, -6.56186e-010, 1.509021e-007, -3.641183e-006,
  1.652839e-009, 9.403711e-012, 4.054786e-008, -9.86068e-007,
  -1.119173e-008, -1.056766e-009, 1.014731e-007, -3.039275e-006,
  1.985346e-009, -9.170444e-011, 2.632317e-008, -8.395209e-007,
  -7.991931e-010, -1.126859e-009, 3.883634e-008, -1.658387e-006,
  2.423743e-009, -8.844915e-011, 1.514645e-008, -5.766502e-007,
  3.193883e-009, -4.611212e-010, 1.128883e-008, -6.499627e-007,
  1.907106e-009, -3.174457e-011, 8.463475e-009, -3.778857e-007,
  1.999946e-009, -1.039354e-010, 2.940956e-009, -2.549147e-007,
  1.34151e-009, -4.075079e-012, 3.605963e-009, -2.465096e-007,
  9.965726e-010, -1.961502e-011, 4.906087e-010, -1.019129e-007,
  9.090859e-010, -3.150239e-012, 1.061674e-009, -1.617104e-007,
  4.918567e-010, -1.70447e-011, 1.624131e-010, -3.595093e-008,
  6.130882e-010, -1.006683e-011, 3.312286e-010, -1.061348e-007,
  2.447781e-010, -1.774359e-011, 2.501249e-010, -6.469129e-009,
  4.191653e-010, -1.647845e-011, 1.667231e-010, -6.978456e-008,
  1.201519e-010, -1.774148e-011, 5.026055e-010, 6.538255e-009,
  2.896212e-010, -2.027279e-011, 3.059305e-010, -4.558464e-008,
  5.53032e-011, -1.258831e-011, 5.259922e-010, 1.15939e-008,
  2.01869e-010, -1.622331e-011, 5.04898e-010, -2.900773e-008,
  2.214941e-011, -6.783487e-012, 4.164738e-010, 1.28602e-008,
  1.412812e-010, -1.070741e-011, 5.049243e-010, -1.794014e-008,
  5.505065e-012, -2.735649e-012, 2.66015e-010, 1.234329e-008,
  9.923675e-011, -5.568334e-012, 4.645081e-010, -1.041211e-008,
  -2.075769e-012, -1.698442e-012, 2.437019e-010, 1.096663e-008,
  6.917423e-011, -4.311987e-012, 5.184145e-010, -5.319353e-009,
  -6.505193e-012, -9.141066e-013, 2.030121e-010, 9.285593e-009,
  4.925578e-011, -3.195831e-012, 5.133862e-010, -2.043112e-009,
  -6.941672e-012, -5.685761e-013, 1.229179e-010, 7.540302e-009,
  3.485523e-011, -2.672059e-012, 4.729078e-010, 3.473165e-011,
  -6.185996e-012, -3.724295e-013, 6.143278e-011, 5.987784e-009,
  2.473072e-011, -1.835588e-012, 3.854588e-010, 1.320427e-009,
  -5.008732e-012, -2.572497e-013, 5.478215e-012, 4.693507e-009,
  1.763573e-011, -8.27332e-013, 2.318356e-010, 2.073736e-009,
  -3.65376e-012, -1.498539e-013, -3.146688e-011, 3.595906e-009,
  1.267126e-011, -7.303328e-016, 7.291618e-011, 2.42741e-009,
  -2.414521e-012, -1.47809e-013, -6.200161e-011, 2.617996e-009,
  9.210446e-012, -1.90208e-014, 9.076416e-011, 2.589065e-009,
  -1.357813e-012, -1.465702e-013, -3.584731e-011, 1.874773e-009,
  6.819205e-012, -1.571815e-013, 8.875502e-011, 2.497021e-009,
  -5.255625e-013, -9.604397e-014, -3.829004e-011, 1.254264e-009,
  5.18125e-012, -1.832112e-013, 1.73098e-011, 2.280936e-009,
  6.585802e-014, -1.905697e-013, -9.452591e-011, 7.550106e-010,
  4.059512e-012, -1.097361e-013, 5.971023e-011, 2.202384e-009,
  5.746309e-013, 2.621116e-014, 4.529117e-011, 6.369253e-010,
  3.301029e-012, -2.803443e-014, 2.434136e-012, 1.929113e-009,
  9.088847e-013, -4.917866e-015, -3.084706e-011, 2.635933e-010,
  2.67573e-012, -7.944403e-014, -2.46723e-011, 1.641641e-009,
  1.109979e-012, -2.916792e-014, -5.112818e-011, 4.482326e-011,
  2.383045e-012, -9.725937e-014, 5.896007e-012, 1.489224e-009,
  1.239774e-012, -2.752266e-014, 1.118501e-011, 3.033548e-011,
  2.132222e-012, 2.134194e-014, 2.269067e-011, 1.338132e-009,
  1.295608e-012, -2.887498e-015, -4.315775e-012, -1.027671e-010,
  1.927665e-012, -1.372745e-014, -2.162909e-011, 1.107755e-009,
  1.306938e-012, 1.905261e-014, 1.771453e-011, -1.096259e-010,
  1.786463e-012, 2.445012e-014, -1.81723e-011, 9.522102e-010,
  1.273257e-012, 3.788009e-014, 2.148491e-013, -1.580014e-010,
  1.658107e-012, -2.816439e-014, -3.734504e-011, 7.801896e-010,
  1.220788e-012, -1.709556e-014, -1.17042e-011, -1.774285e-010,
  1.554036e-012, -1.873781e-014, -2.418014e-012, 7.230113e-010,
  1.145923e-012, -2.678563e-014, -2.416637e-011, -2.081229e-010,
  1.468902e-012, -4.205094e-014, 7.356587e-013, 6.188602e-010,
  1.068955e-012, -2.86004e-014, -3.244988e-011, -2.17357e-010,
  1.384848e-012, -1.001463e-014, 7.454236e-012, 5.375891e-010,
  9.960396e-013, 4.510846e-015, 5.96411e-012, -1.535776e-010,
  1.304212e-012, 4.715706e-014, -4.343341e-012, 4.767686e-010,
  9.148127e-013, 3.457893e-014, 1.279981e-011, -1.32938e-010,
  1.229515e-012, 5.468362e-014, -2.234376e-011, 3.935406e-010,
  8.388222e-013, 4.253857e-014, 6.003934e-012, -1.308517e-010,
  1.154887e-012, 3.679729e-014, -1.584204e-011, 3.522121e-010,
  7.579219e-013, 3.683513e-014, -7.30246e-012, -1.326446e-010,
  1.102645e-012, 4.074695e-014, -1.612705e-011, 2.94407e-010,
  7.005517e-013, -8.561322e-015, -2.080108e-011, -1.295244e-010,
  1.013304e-012, -2.613007e-014, 1.506557e-012, 2.799953e-010,
  6.304489e-013, -6.26277e-014, -4.757338e-011, -1.377303e-010,
  9.389498e-013, -8.796527e-014, 4.44658e-011, 2.994129e-010,
  5.528633e-013, -1.378514e-013, -2.21861e-011, -1.083846e-010,
  8.760528e-013, -8.09747e-014, 6.990606e-011, 3.342995e-010,
  5.686319e-013, 2.290764e-013, 1.044799e-010, 1.094242e-010,
  8.303193e-013, 4.746622e-014, 2.985589e-011, 2.458108e-010,
  3.471594e-013, -2.624823e-014, -2.51121e-011, -1.143114e-010,
  7.245897e-013, -1.050237e-013, 2.969491e-012, 1.733243e-010,
  4.154771e-013, -9.462341e-014, -4.40586e-012, -5.346376e-011,
  6.888685e-013, -1.622007e-013, 5.021495e-011, 2.331655e-010,
  3.958712e-013, -7.481125e-014, -1.486561e-011, -9.497136e-011,
  6.328833e-013, -1.434172e-013, 5.333949e-012, 1.617313e-010,
  3.774483e-013, -2.545659e-014, 4.683032e-011, 3.148163e-011,
  6.306351e-013, 4.078207e-014, 2.437094e-011, 1.886432e-010,
  3.73536e-013, 1.801445e-014, 3.714429e-011, 3.204448e-011,
  6.576555e-013, 2.052825e-014, -1.580055e-011, 1.161113e-010,
  3.438815e-013, 5.792836e-014, 1.358363e-011, -1.489836e-011,
  5.617792e-013, -1.976757e-014, -4.979741e-011, 4.65975e-011,
  3.046354e-013, -1.771063e-014, -3.274608e-012, -3.110519e-011,
  5.194072e-013, -3.577034e-014, -3.474875e-012, 1.047169e-010,
  2.804722e-013, -1.96676e-014, -3.37067e-012, -3.88833e-011,
  4.814528e-013, -5.514346e-014, 3.820471e-011, 1.732206e-010,
  2.761257e-013, -8.595186e-014, -4.611266e-011, -9.577372e-011,
  4.004408e-013, -6.97003e-014, 3.338608e-011, 1.67449e-010,
  2.49396e-013, -6.880525e-014, -9.726327e-012, -3.261223e-011,
  3.915958e-013, -4.676183e-014, 2.959451e-011, 1.417035e-010,
  2.356119e-013, -2.563051e-015, 8.090723e-011, 1.154466e-010,
  3.98721e-013, 4.964803e-014, 9.736465e-012, 9.208721e-011,
  2.305267e-013, -2.755469e-014, -1.73506e-012, -1.678016e-011,
  3.709067e-013, -3.28395e-014, -1.853469e-012, 7.250137e-011,
  2.03358e-013, -3.320412e-014, 1.816228e-011, 2.602285e-011,
  3.562652e-013, -5.378101e-014, 1.978053e-011, 9.840765e-011,
  2.176325e-013, -4.204032e-014, -2.557623e-011, -4.476024e-011,
  3.716732e-013, -3.498937e-014, -7.905309e-013, 5.026277e-011,
  1.946587e-013, 2.70415e-014, 1.134204e-010, 1.773737e-010,
  3.321568e-013, 7.282424e-014, -1.753841e-011, 1.463044e-011,
  1.839765e-013, 4.536653e-014, 4.929581e-011, 8.062622e-011,
  3.048936e-013, 2.944471e-014, -8.342273e-012, 4.415089e-011,
  1.450308e-013, -1.784463e-013, -3.126478e-012, -2.366875e-011,
  2.871087e-013, -3.728639e-014, 8.256882e-011, 2.272642e-010,
  2.312741e-013, -4.263447e-014, -1.13729e-011, -4.713693e-011,
  3.705252e-013, -8.122433e-014, 2.541678e-011, 9.812742e-011,
  1.456133e-013, -6.35358e-015, -3.078952e-011, -6.128665e-011,
  2.439968e-013, -1.053417e-013, -3.195473e-011, -1.918557e-011,
  1.407006e-013, -3.324249e-014, 5.682582e-011, 1.0989e-010,
  2.56438e-013, 6.121653e-014, 4.643273e-011, 9.756462e-011,
  1.54529e-013, 5.517487e-014, 1.475482e-010, 2.297266e-010,
  2.58166e-013, 1.686799e-013, 6.233355e-011, 1.358018e-010,
  1.737623e-013, -3.690243e-014, 6.763222e-012, -9.246187e-012,
  1.550166e-013, -5.343692e-014, 6.839916e-012, 3.39401e-011,
  1.239358e-013, -6.096556e-014, 7.706808e-012, 7.360732e-012,
  2.031784e-013, -6.883737e-014, 4.834771e-011, 9.784181e-011,
  1.173318e-013, -3.723959e-014, -3.19531e-011, -6.993353e-011,
  1.78793e-013, -1.262957e-013, 1.188826e-011, 4.344974e-011,
  1.012847e-013, -2.187979e-014, 5.249572e-012, -4.096876e-012,
  1.848769e-013, -5.934143e-014, 1.28959e-011, 2.942036e-011,
  4.799176e-014, -1.877239e-014, -3.241388e-013, -5.477062e-012,
  2.074823e-013, -4.375063e-014, 1.178609e-011, 4.465236e-011,
  8.314252e-014, -9.10926e-015, 2.240828e-012, -1.003877e-011,
  1.815024e-013, -3.994203e-014, -2.46254e-012, 2.522182e-011,
  1.010668e-013, -3.051623e-014, 4.554381e-012, -5.885033e-012,
  1.622167e-013, -2.493198e-014, 5.407561e-013, 3.2698e-011,
  9.626851e-014, -2.571131e-014, -6.673531e-012, -2.254208e-011,
  1.512069e-013, -4.096499e-014, 1.380859e-012, 3.700625e-011,
  8.934548e-014, -4.608504e-014, -1.257796e-011, -3.355036e-011,
  1.507598e-013, -4.024484e-014, 2.511176e-011, 6.161922e-011,
  9.172371e-014, -9.86801e-015, 2.865112e-011, 6.335613e-011,
  1.509971e-013, 1.429147e-014, 3.296745e-012, 2.359891e-011,
  8.561381e-014, -1.108485e-014, -2.139536e-011, -3.707629e-011,
  1.292226e-013, -5.906252e-014, -1.042409e-011, 2.279093e-011,
  8.199265e-014, 1.797428e-015, -2.189346e-011, -4.543408e-011,
  1.215482e-013, -7.102695e-014, -3.741397e-011, -3.364197e-011,
  9.121705e-014, -4.007039e-014, -2.622165e-011, -4.511103e-011,
  1.066536e-013, -1.416211e-014, 3.307323e-012, 3.577996e-011,
  1.088625e-013, 1.50765e-014, 9.745452e-012, 2.537806e-011,
  6.472981e-015, 1.780291e-014, -5.53782e-011, -7.753417e-011,
  8.427263e-014, 9.055775e-014, 3.159781e-011, 5.286144e-011,
  1.182364e-013, -5.854131e-015, -4.641437e-011, -6.146115e-011,
  8.86961e-014, 3.846116e-014, -1.153455e-010, -2.002644e-010,
  9.133933e-014, -8.09548e-014, -5.4876e-012, 3.229083e-011,
  1.076901e-013, -1.858994e-014, -1.53598e-010, -2.520956e-010,
  1.189772e-013, -1.072212e-013, 2.620866e-012, 3.353198e-011,
  -3.277003e-014, -1.002033e-013, -3.868517e-011, -7.940514e-011,
  1.298393e-013, 1.438779e-014, 6.62404e-011, 9.274478e-011,
  4.786134e-014, 4.474664e-014, 4.207435e-011, 8.941786e-011,
  8.857289e-014, -6.636004e-014, -1.666201e-012, 4.233712e-012,
  2.616829e-014, -3.523345e-013, 3.79975e-011, 4.371236e-011,
  1.928771e-013, -1.136596e-013, 7.183341e-011, 8.575855e-011,
  9.122781e-014, -2.117037e-014, -2.957735e-011, -3.070094e-011,
  1.075786e-013, 1.044459e-014, 2.916981e-011, 7.514346e-011,
  1.043215e-013, -2.192677e-014, 8.499114e-012, 3.361086e-011,
  1.714375e-013, -5.224364e-014, 4.24862e-011, 1.213079e-010,
  2.233426e-014, -3.04054e-014, 2.522629e-012, 2.545052e-011,
  8.752417e-014, -2.439099e-014, -2.323269e-011, -3.882931e-011,
  -5.035368e-015, -4.742314e-014, -6.611005e-011, -3.172962e-011,
  9.027058e-015, 1.744392e-014, 5.532876e-011, 8.682521e-011,
  -2.607069e-014, -6.104894e-014, -7.104301e-011, -1.208094e-010,
  5.304748e-014, -3.916515e-014, 3.852084e-011, 4.986475e-011,
  -8.632622e-014, -1.563771e-013, 4.121163e-011, 9.992408e-011,
  1.692784e-013, -5.941539e-014, 3.08205e-011, 3.627307e-011,
  1.340621e-013, -2.034684e-014, -5.155461e-011, -1.200133e-010,
  2.112988e-013, -1.623528e-015, 7.41334e-011, 1.226302e-010,
  4.644732e-014, 7.317149e-016, 8.77141e-011, 2.141393e-010,
  -1.21798e-013, 3.451687e-014, 3.817049e-011, 1.098783e-010,
  9.477683e-014, 3.418773e-014, 4.600234e-011, 4.445451e-011,
  1.328571e-013, -3.8493e-016, -3.27876e-011, -1.87633e-011,
  2.23455e-014, -1.258559e-014, 4.108007e-011, 8.596501e-011,
  5.369576e-014, 2.81804e-014, 2.047993e-011, 2.791136e-011,
  1.260916e-013, -1.088484e-014, -3.731683e-012, 7.801134e-012,
  -1.152458e-014, 2.229344e-014, 5.296476e-011, 1.143939e-010,
  -1.01141e-013, -2.45713e-014, -6.71697e-011, -9.212846e-011,
  1.13641e-013, -8.972597e-014, 2.119558e-011, -2.551328e-012,
  1.433799e-014, -2.764727e-014, -8.638551e-012, -5.165752e-012,
  6.810854e-014, -1.890768e-014, -2.247346e-012, 1.415773e-011,
  3.543257e-014, -1.209389e-014, 8.121326e-012, 1.253661e-011,
  5.779814e-014, 4.267213e-015, 2.056064e-011, 4.343327e-011,
  1.299363e-013, 4.474602e-015, -3.542905e-011, -6.655139e-011,
  8.436042e-014, -1.60428e-014, -1.649854e-011, -1.179616e-011,
  2.441074e-014, -2.335219e-014, -1.391076e-011, -2.201758e-011,
  5.037372e-014, -3.036493e-014, 1.886649e-011, 3.489019e-011,
  3.801639e-014, -5.504778e-015, 1.679968e-012, -8.351665e-012,
  4.609022e-014, -7.238081e-015, -1.166326e-011, -2.164548e-011,
  3.46335e-014, -1.331942e-014, -4.517962e-012, -1.322163e-011,
  4.637743e-014, -1.40673e-014, -1.869467e-011, -2.488765e-011,
  2.701971e-014, -1.525799e-014, -1.035869e-011, -1.796683e-011,
  5.248617e-014, -1.800355e-014, 5.821354e-012, 1.75551e-011,
  2.678792e-014, -9.44821e-015, -5.752585e-012, -8.245332e-012,
  4.784149e-014, -1.533481e-014, -1.652584e-012, 5.144848e-012,
  2.997872e-014, -1.698739e-014, -2.537074e-012, -7.036588e-012,
  4.823503e-014, -2.473084e-014, 6.8623e-012, 1.317137e-011,
  1.870611e-014, -2.49271e-014, -1.14468e-011, -1.766716e-011,
  5.579903e-014, -2.878141e-014, 1.85742e-011, 2.165107e-011,
  2.115497e-015, -1.681466e-014, 3.533071e-012, -2.408829e-012,
  7.078207e-016, -2.007808e-014, -3.265537e-013, 3.982518e-012,
  2.717997e-015, -1.128899e-014, 6.271792e-012, 1.227005e-011,
  3.02584e-014, -2.229102e-014, -8.617686e-013, -1.295856e-011,
  4.396036e-014, 6.822718e-014, 1.877205e-012, -7.797265e-012,
  5.615452e-014, -3.781295e-014, -6.464741e-011, -1.206545e-010,
  4.365048e-014, 1.5052e-014, 1.138948e-011, 2.214407e-011,
  4.604403e-014, 2.067336e-015, 1.698896e-011, 2.040937e-011,
  1.319721e-014, -6.157708e-015, 5.693793e-012, 5.323474e-012,
  6.744744e-014, -1.754772e-014, 1.334702e-011, 1.796612e-011,
  3.540752e-014, 3.699633e-014, 1.744909e-011, 2.723158e-011,
  9.132294e-014, -3.318899e-014, -1.019051e-011, -3.601203e-011,
  1.206344e-014, -1.83241e-014, 9.367301e-012, 3.538724e-011,
  7.266178e-016, 6.573291e-015, 3.55171e-011, 6.655001e-011,
  -1.047128e-013, -1.053352e-014, 6.659456e-011, 1.094895e-010,
  2.900092e-014, 9.50723e-016, 3.215169e-011, 1.694978e-012,
  6.544401e-014, -6.210828e-015, -9.072497e-012, -1.619585e-011,
  4.343259e-014, -4.8845e-015, -4.063046e-012, 1.932655e-011,
  8.867265e-014, -1.530288e-014, 8.317797e-011, 9.456581e-011,
  -5.64757e-014, 9.418257e-015, -2.391035e-011, -5.639803e-011,
  -1.720619e-013, 2.514133e-014, 1.571422e-012, 1.912945e-011,
  3.744976e-014, -1.455434e-014, -5.510797e-011, -1.283004e-010,
  -8.322357e-015, 5.905359e-015, -4.573482e-011, -5.26775e-011,
  -9.288437e-015, 1.304999e-015, -5.097382e-011, -7.731663e-011,
  9.481908e-014, 2.07097e-014, -1.252246e-011, 4.304075e-011,
  -2.214765e-013, 3.420539e-014, -2.482889e-011, 2.870535e-011,
  2.890348e-013, -3.836129e-014, 2.202211e-011, 3.800249e-011,
  8.206311e-014, -2.260648e-014, 5.058899e-011, 1.245991e-010,
  1.658799e-014, 7.944251e-016, 7.71557e-011, 1.388574e-010,
  1.012533e-013, -2.580801e-014, -6.012518e-011, -9.49241e-011,
  7.521189e-014, 1.155778e-014, 6.235978e-011, 1.142919e-010,
  4.076121e-014, 2.471681e-014, -5.760925e-011, -9.42868e-011,
  1.772003e-013, -4.776775e-015, 3.796504e-011, 1.954827e-011,
  3.183617e-014, 2.478559e-015, -1.148442e-010, -1.322358e-010,
  -4.244666e-014, 9.070664e-014, 2.051102e-011, 2.307706e-011,
  3.020093e-015, -1.315098e-013, -1.881102e-010, -3.730834e-010,
  -1.109142e-013, -1.276357e-013, 4.493531e-011, 3.717456e-011,
  1.141639e-013, 6.866618e-014, 4.507668e-011, 9.170497e-011,
  1.133657e-013, -3.897719e-015, -6.787729e-011, -1.555471e-010,
  6.973185e-014, -1.026929e-013, -1.145397e-010, -1.455801e-010,
  -9.948615e-014, -6.430245e-015, -2.29045e-011, 1.146647e-011,
  -1.479731e-013, -1.996485e-013, -9.563636e-011, -1.405214e-010,
  -1.454582e-013, -3.673615e-014, -1.719262e-011, 2.693279e-011,
  4.583137e-013, 1.193767e-014, 2.597049e-011, -5.400546e-011,
  1.9043e-014, -7.891849e-014, -1.144558e-010, -1.835015e-010,
  -8.344363e-014, -9.520797e-015, 1.516596e-010, 2.212093e-010,
  1.395306e-014, 2.818605e-014, 6.526979e-012, 3.193427e-012,
  3.140672e-014, 2.186239e-014, 2.457455e-011, 3.293511e-011,
  -8.27809e-015, 9.178018e-015, 3.935238e-012, 1.773424e-011,
  1.085876e-014, 1.623682e-014, 2.041164e-011, 3.099666e-011,
  1.022052e-013, 1.542845e-014, -1.186428e-011, -4.229288e-011,
  7.689061e-014, -1.27596e-014, -2.140565e-012, 9.383066e-012,
  6.775693e-014, -1.648219e-015, 2.357378e-011, 4.883273e-011,
  -3.738522e-014, 4.323353e-015, -6.620115e-012, -2.327527e-011,
  6.522508e-015, 1.683169e-014, 1.067289e-011, 2.598975e-011,
  -1.248238e-014, 1.124644e-014, 2.084543e-011, 1.546914e-011,
  4.355264e-014, -2.527489e-015, 1.65703e-011, 2.690766e-011,
  2.024244e-014, -2.873288e-015, 4.470795e-012, 4.970054e-012,
  4.167789e-014, -1.885785e-014, 3.238015e-011, 4.940138e-011,
  3.35271e-014, -8.347463e-016, -1.150731e-011, -8.711656e-012,
  -5.202037e-014, 5.470206e-015, -1.474869e-011, -9.986174e-012,
  3.264131e-014, -4.178561e-015, -1.842897e-011, -1.710877e-011,
  -1.098454e-015, 1.24802e-014, -1.425098e-011, -2.746516e-011,
  2.511304e-014, -3.83086e-014, 2.385319e-012, -7.466064e-012,
  -5.349842e-014, -2.829681e-014, 4.94723e-011, 9.935111e-011,
  -9.815815e-015, 2.267956e-014, -1.396402e-011, -4.154524e-011,
  -1.138253e-013, -5.814841e-014, -3.347205e-011, -6.708786e-011,
  4.534771e-014, 8.131389e-014, -2.339338e-011, -8.08243e-012,
  1.060183e-014, 1.57361e-014, 1.853118e-011, 4.748804e-012,
  5.95761e-014, -7.633602e-014, 1.315748e-011, 2.496279e-011,
  1.903124e-014, -2.753015e-014, 2.034494e-011, 1.990512e-011,
  6.693033e-014, -6.343657e-015, -9.924029e-013, 6.332197e-012,
  3.669435e-014, 3.364904e-015, -4.814529e-012, -2.820954e-011,
  4.404382e-014, -4.675055e-014, -1.199008e-011, -1.94341e-011,
  8.804073e-014, -5.196874e-014, -5.51513e-011, -1.036834e-010,
  4.149311e-014, 4.676006e-014, 4.118273e-011, 1.044851e-010,
  -1.370134e-013, 3.381749e-015, -1.562681e-011, -6.299592e-011,
  4.197862e-014, -1.09375e-014, 2.82793e-011, 3.9648e-011,
  5.048058e-014, 1.910825e-014, 3.826389e-011, 2.193595e-011,
  9.937206e-014, -9.703584e-015, -1.416292e-011, 1.220247e-011,
  2.109311e-014, -4.232283e-015, -9.757451e-012, -3.631611e-011,
  9.229005e-014, -2.716792e-014, -6.206823e-011, -9.11159e-011,
  6.893911e-015, -5.35447e-014, 1.118117e-011, 2.474609e-011,
  5.160379e-014, -8.087463e-015, 1.467579e-011, 5.610837e-011,
  5.753188e-014, -1.500971e-014, 3.354825e-011, 2.810315e-011,
  8.533456e-014, -1.202037e-014, 2.857256e-011, 4.939419e-011,
  -1.49369e-013, 1.291907e-014, 3.103756e-011, 1.204671e-010,
  -1.428815e-013, -9.41385e-015, -5.138396e-011, -8.80677e-011,
  1.027404e-014, 3.257689e-014, 3.825014e-011, 1.132139e-010,
  1.66029e-014, 3.245944e-014, 1.043172e-011, 8.388309e-012,
  7.970781e-015, -4.187338e-015, -3.520393e-011, -5.869981e-011,
  8.315402e-014, -3.417337e-014, -6.343426e-011, -8.321138e-011,
  -9.353593e-015, 2.630785e-014, -7.441448e-012, 1.95745e-011,
  -5.874684e-014, -1.186994e-014, -2.222683e-011, -3.373277e-011,
  5.752971e-014, -1.565875e-014, -6.119843e-012, 8.630297e-012,
  4.785419e-014, -1.504895e-014, 2.902409e-012, 4.081802e-013,
  3.246243e-015, -7.457259e-015, -2.604406e-011, -5.502852e-011,
  2.386551e-014, -2.527171e-014, -1.092641e-012, -1.504129e-011,
  -2.587902e-014, 7.071356e-016, -1.036381e-011, -2.031995e-011,
  1.620069e-014, -5.314384e-014, -3.803854e-011, -5.842259e-011,
  -8.912954e-014, -2.272774e-014, -2.451111e-011, -6.665898e-011,
  9.695189e-014, 3.776972e-016, -1.529312e-011, -7.788951e-011,
  -1.16611e-014, -1.512834e-014, 2.073092e-011, -5.067166e-012,
  1.675862e-015, -3.441365e-014, -3.544796e-011, -4.935795e-011,
  6.298115e-015, -3.840336e-014, 1.274698e-011, 2.497216e-011,
  -8.588878e-015, -1.652811e-014, -1.676116e-012, 3.225354e-011,
  -3.555719e-014, -5.244121e-014, -9.054469e-013, 2.440717e-013,
  5.799252e-014, -1.888125e-014, 9.576199e-013, -7.285953e-012,
  2.692955e-014, 6.982549e-015, 3.953144e-011, 5.767617e-011,
  -1.595509e-014, 4.915961e-014, 6.423177e-012, 3.538887e-011,
  4.07011e-014, -1.651488e-014, 3.050512e-011, 3.831305e-011,
  -4.135891e-014, 2.194423e-014, -1.089948e-011, -5.832438e-012,
  -5.516018e-015, -5.056006e-014, -1.933319e-011, -1.734432e-011,
  8.743821e-014, -9.478519e-015, 2.965155e-011, 6.09413e-011,
  1.772094e-013, 5.534305e-014, 3.152387e-011, 8.387754e-011,
  -9.556022e-014, 4.710966e-015, 6.550111e-011, 1.876318e-010,
  2.226845e-013, -5.110174e-014, 5.493035e-011, 1.217287e-010,
  -2.70334e-013, -8.620606e-014, 4.38856e-011, 2.166851e-010,
  1.381383e-013, -6.20006e-014, 5.686356e-011, 8.164961e-011,
  -1.578038e-013, 5.455623e-014, 2.032861e-012, 9.026018e-011,
  2.59552e-013, 2.408707e-014, 1.60393e-010, 2.149118e-010,
  -6.76106e-014, 4.400826e-014, 3.816196e-011, 1.179073e-010,
  -1.713668e-013, 5.360182e-014, 7.89204e-011, 1.538887e-010,
  -7.151471e-014, 9.605649e-015, 4.302287e-011, 1.959564e-011,
  8.176269e-014, 3.723711e-015, 1.980425e-011, 3.310837e-011,
  3.464908e-014, -1.30022e-014, -2.751668e-011, -4.390836e-011,
  1.480048e-014, -2.302773e-015, 5.637509e-011, 9.810801e-011,
  -6.093193e-014, -4.769089e-014, 1.634651e-011, 6.952933e-011,
  1.420708e-013, -2.142769e-014, -6.437498e-011, -1.705508e-010,
  5.247733e-014, -5.673665e-014, 1.130952e-010, 2.34284e-010,
  8.388632e-014, -3.000586e-014, 7.795136e-011, 1.596219e-010,
  -8.958096e-014, 3.484169e-014, 4.484405e-011, 1.076953e-010,
  8.36642e-014, -6.336172e-015, 9.332377e-012, 8.265959e-011,
  -8.839583e-014, 4.555263e-015, -3.546214e-011, -3.302025e-011,
  1.695836e-014, 1.804669e-014, 2.789722e-011, -1.264631e-011,
  6.95346e-014, -1.584345e-014, -3.868632e-011, -5.02785e-011,
  1.43714e-013, -6.491548e-014, -4.701896e-012, -2.038771e-011,
  -3.360759e-014, -9.207725e-016, 8.750184e-011, 1.987066e-010,
  -1.528754e-014, 2.056249e-014, -1.044761e-011, -2.008116e-011,
  2.509592e-014, -3.013451e-014, -3.91718e-011, -4.091672e-011,
  -6.466647e-014, -2.155527e-014, 2.329428e-011, 3.981856e-011,
  1.455188e-015, 3.57668e-015, 3.584606e-011, 5.534926e-011,
  -1.016923e-014, 5.454478e-014, 2.754371e-012, 4.588463e-012,
  4.49277e-014, -1.029775e-014, -6.466749e-011, -1.287025e-010,
  -1.340543e-013, 4.695094e-014, 2.812684e-011, 6.073855e-011,
  1.156801e-013, -1.496553e-014, -5.745476e-011, -9.610695e-011,
  1.883424e-014, -4.492557e-015, 5.18218e-011, 7.620843e-011,
  4.717873e-014, 1.244511e-015, 1.698655e-011, 2.741085e-011,
  -2.214379e-014, -1.747242e-014, 3.516125e-011, 9.384619e-011,
  -7.462238e-014, 1.987733e-014, 6.936862e-011, 1.145057e-010,
  -8.150403e-014, 2.861074e-014, 1.070452e-010, 3.038457e-010,
  -2.964488e-013, 3.67765e-014, -4.030959e-011, -7.839842e-011,
  -1.291216e-013, -2.929757e-014, 1.124425e-011, -1.336181e-012,
  -2.213124e-014, 6.175742e-015, -2.682922e-011, -6.309429e-011,
  -4.849819e-014, -2.030812e-014, 1.626565e-011, -1.556282e-011,
  2.758074e-014, 1.725557e-014, -1.691351e-011, -3.32312e-011,
  -7.879782e-014, -6.654475e-015, 9.118619e-011, 1.292929e-010,
  1.903499e-013, -4.442183e-014, -6.944627e-011, -1.406694e-010,
  2.492698e-014, -7.894219e-014, -2.747612e-010, -5.868386e-010,
  5.581858e-013, -5.237915e-014, 3.985342e-012, -2.065476e-010,
  3.580115e-014, -1.070717e-014, -1.443106e-010, -2.394607e-010,
  -9.837413e-014, -8.021183e-014, -4.379399e-012, -1.910915e-011,
  -2.595933e-013, 2.171136e-015, -1.907328e-011, 2.48553e-011,
  -2.012424e-013, 5.847054e-014, 8.817975e-011, 8.449048e-011,
  7.777066e-015, 1.38163e-013, 1.238303e-010, 3.49059e-010,
  -1.099166e-013, -9.19358e-014, -6.829839e-011, -9.479497e-011,
  -1.181639e-013, -1.222743e-014, -9.000774e-011, -1.14666e-010,
  6.264038e-014, -5.153649e-014, -2.211552e-011, -9.643661e-011,
  5.379843e-014, -2.292858e-014, -4.44378e-011, -5.369182e-011,
  5.085419e-014, -6.168895e-014, -6.205001e-012, -4.460002e-011,
  1.434564e-014, 1.296037e-015, 2.422501e-012, -2.816929e-013,
  1.8545e-014, 4.376407e-015, -1.665522e-012, 4.765327e-012,
  4.248274e-014, -3.781232e-015, 4.749964e-011, 2.461277e-011,
  -4.523727e-015, 5.527519e-015, -2.426964e-011, -3.915923e-012,
  6.513174e-014, -5.64814e-015, -8.339955e-012, -5.762543e-012,
  -6.962721e-014, 1.526343e-014, 1.091623e-011, 1.379251e-011,
  9.121927e-015, -4.915019e-015, -4.575864e-012, -9.898947e-012,
  2.261623e-014, -5.0982e-015, 3.945887e-012, 1.329919e-011,
  1.134771e-014, 5.267246e-016, -5.10419e-012, -1.029871e-011,
  1.94438e-014, -1.772395e-015, -7.748658e-012, 3.427367e-012,
  1.477198e-014, 3.54235e-015, -1.412108e-011, -7.974827e-012,
  2.285159e-014, -6.136262e-016, -4.326507e-013, -4.546086e-012,
  5.29585e-014, -3.051362e-016, -6.07641e-012, -8.480236e-012,
  9.518297e-014, -1.518201e-014, -9.269174e-012, -1.430119e-012,
  1.091068e-014, -2.047589e-016, -1.17001e-011, -1.745781e-011,
  1.755289e-014, -5.757054e-015, 1.033264e-012, 9.688669e-012,
  1.730798e-014, 6.076058e-015, 8.166936e-012, -3.822842e-012,
  2.453262e-014, 1.130012e-015, 9.231923e-012, -1.765584e-012,
  8.950475e-015, -7.638354e-014, 1.555781e-011, 5.47768e-013,
  3.068373e-014, 3.817436e-014, 1.981837e-011, 7.11847e-012,
  9.814033e-014, -1.256364e-014, -1.758589e-013, 1.516856e-012,
  3.437778e-015, -6.087402e-015, -2.332298e-012, 3.150029e-012,
  2.163649e-014, -1.101677e-015, 1.987163e-012, -2.121895e-013,
  2.128545e-014, 1.452586e-015, -3.456901e-012, 2.792536e-012,
  1.821394e-014, 2.003605e-015, -2.902027e-012, -5.925606e-012,
  2.712585e-014, 3.104805e-015, -3.397349e-012, 8.54343e-012,
  1.605862e-014, -4.412552e-016, 1.204106e-012, -1.919753e-012,
  2.646183e-014, 7.059465e-015, -4.747653e-012, 4.921734e-012,
  1.525374e-014, 8.019699e-016, 2.778896e-012, 1.065718e-012,
  2.948378e-014, 3.701895e-015, 1.587717e-012, 8.513914e-012,
  2.008623e-014, -1.650055e-015, -2.492505e-012, -3.536163e-012,
  3.163279e-014, 1.854735e-015, 9.235964e-013, 8.951009e-012,
  2.630943e-014, 1.422512e-015, 8.430781e-014, -4.760536e-012,
  2.511449e-014, 2.377531e-015, -6.122245e-014, 1.021708e-011,
  1.540159e-014, 2.762241e-015, 2.885528e-013, -2.895004e-012,
  2.519903e-014, 5.621873e-015, -1.279439e-012, 4.955371e-012,
  1.615873e-014, -2.702582e-015, 1.914569e-012, -6.76824e-014,
  2.914719e-014, 7.567746e-015, 2.105443e-013, 7.251153e-012,
  2.015433e-014, -2.270875e-015, 9.687083e-013, 6.763841e-013,
  3.377427e-014, 4.26099e-015, -6.1309e-012, -1.03105e-013,
  2.006527e-014, -4.319387e-017, -1.067384e-013, -8.945979e-013,
  3.112089e-014, 1.546315e-015, 2.857142e-012, 9.868026e-012,
  2.175951e-014, 2.162987e-015, -3.824855e-012, -1.979072e-012,
  3.120151e-014, -1.551098e-015, 8.205523e-012, 1.632103e-011,
  3.313996e-014, 5.296723e-016, -8.665315e-012, -6.278571e-012,
  2.410444e-014, -1.374444e-016, 6.366998e-012, 2.118783e-011,
  8.136822e-014, -9.567433e-015, 2.710846e-012, -6.281683e-013,
  -1.135299e-014, 6.543853e-015, -2.020298e-012, 4.875454e-012,
  2.449107e-014, 3.235212e-015, -5.962333e-012, -4.61135e-012,
  3.228433e-014, -1.516168e-014, 3.84627e-012, 9.898458e-012,
  2.297803e-014, 2.564508e-015, 1.329631e-011, 7.824325e-012,
  4.13017e-014, -5.170919e-015, -9.582705e-012, 3.026993e-012,
  2.270434e-014, 8.660288e-015, 9.647292e-012, 9.021141e-012,
  4.278687e-014, -1.175741e-014, -4.801679e-012, 7.585202e-012,
  1.813692e-015, 1.43299e-015, -5.72492e-012, -3.960898e-012,
  -5.460437e-014, 1.219189e-014, 9.036968e-013, 1.205928e-011,
  2.990675e-014, -3.590454e-017, -3.697396e-012, -2.59235e-012,
  3.691784e-014, -6.100234e-016, 9.13176e-012, 1.544561e-011,
  2.90664e-014, -2.708663e-015, -6.743328e-012, -5.601825e-012,
  3.959915e-014, -6.067021e-015, 1.54195e-011, 1.773864e-011,
  3.641241e-014, -1.665858e-015, -4.290471e-012, -1.40782e-012,
  4.297127e-014, -4.949365e-015, -2.979861e-013, 7.400169e-012,
  2.20913e-014, -1.14796e-015, -2.560809e-012, -4.592465e-011,
  4.324076e-014, -2.246765e-015, -4.003422e-014, 1.425533e-011,
  2.798656e-014, -5.59211e-015, 1.947242e-012, -8.612117e-013,
  3.877636e-014, -9.57047e-016, 2.472571e-012, 1.07043e-011,
  1.455541e-014, -2.00548e-015, 1.479837e-011, 2.930831e-011,
  2.90093e-014, -3.236199e-015, -2.256239e-012, -7.428968e-012,
  2.280535e-014, -1.42768e-016, 8.781737e-012, 1.058807e-011,
  4.561374e-014, -7.672181e-015, -1.420749e-012, -6.759564e-013,
  -5.097864e-015, 1.541586e-015, 1.011306e-012, 3.415579e-012,
  1.177277e-013, -1.830353e-014, -6.222384e-012, 3.377828e-012,
  1.699107e-014, -3.262847e-015, -1.423156e-011, -2.051119e-011,
  1.386818e-013, -1.673187e-014, 3.247355e-012, 1.959902e-011,
  3.176945e-014, -1.303655e-015, -1.178082e-012, -4.465616e-012,
  5.754839e-014, -6.750866e-015, 3.238083e-012, 1.576211e-011,
  3.657352e-014, -2.978776e-016, -1.261997e-012, -4.007464e-012,
  6.083967e-014, -5.968512e-015, 7.43945e-013, 1.390836e-011,
  4.464469e-014, -5.462643e-015, -8.592535e-013, -4.51618e-012,
  7.212023e-014, -3.002166e-015, 1.707787e-013, 1.60664e-011,
  6.864483e-014, -3.628049e-015, -3.719953e-012, -7.549446e-012,
  1.013012e-013, -6.407878e-015, 5.999187e-012, 1.929786e-011,
  3.320289e-014, 1.973344e-015, 2.972028e-012, -2.347447e-012,
  6.132616e-014, -3.582052e-015, 9.945652e-013, 1.331437e-011,
  4.145088e-014, -9.167068e-016, 3.995328e-012, 4.45768e-012,
  6.747708e-014, 2.183879e-015, 2.237123e-012, 1.754699e-011,
  3.994691e-014, 1.988413e-015, 1.05813e-012, -3.586434e-012,
  6.782193e-014, 2.967737e-015, 1.201901e-012, 1.885434e-011,
  1.32339e-013, -9.377169e-015, 2.292286e-013, -3.540184e-012,
  3.207314e-014, 9.868849e-015, 4.186486e-013, 2.079471e-011,
  4.761852e-014, 5.31154e-015, 9.709285e-013, -3.64739e-012,
  7.278207e-014, 2.952696e-015, 1.840461e-012, 2.186755e-011,
  4.227924e-014, -1.297632e-014, -4.109688e-013, -1.749606e-012,
  8.113412e-014, 3.039815e-014, 6.981968e-013, 2.365285e-011,
  4.514465e-014, 1.781727e-015, 1.311815e-012, -4.545035e-012,
  7.665974e-014, 1.160642e-014, -3.008607e-012, 1.573538e-011,
  8.741226e-014, -5.717151e-014, -1.400562e-012, -1.105128e-012,
  2.102619e-013, 1.77654e-014, -1.006633e-011, 2.264703e-011,
  5.98979e-014, 9.330303e-015, -7.990277e-014, 3.059641e-013,
  9.695428e-014, 1.438076e-014, -5.26372e-012, 2.796919e-011,
  5.057772e-014, 7.097511e-015, 2.632424e-012, -7.896179e-012,
  8.574922e-014, 1.754655e-014, -4.301976e-012, 2.235797e-011,
  4.956049e-014, 8.044537e-015, 1.134724e-012, -5.286151e-012,
  8.860287e-014, 1.226783e-014, -6.952883e-013, 2.384266e-011,
  6.157671e-015, 1.403189e-014, -2.753562e-012, -8.529408e-012,
  8.003181e-014, 8.199803e-015, 9.240783e-013, 2.418859e-011,
  2.852408e-014, 1.36104e-014, 2.996566e-012, -1.545265e-012,
  9.818844e-014, 1.57025e-014, -3.515867e-012, 3.233173e-011,
  6.329875e-014, 5.955345e-015, 6.207905e-013, -4.3906e-012,
  9.840892e-014, 9.042259e-015, -4.957413e-012, 2.273187e-011,
  6.078614e-014, 5.323411e-015, -1.953231e-012, -8.492776e-012,
  1.104203e-013, 5.638013e-015, -3.866414e-012, 2.488308e-011,
  5.842677e-014, 7.730019e-015, -1.203836e-012, -7.142445e-012,
  1.344483e-013, -1.209995e-015, 3.957341e-012, 3.423025e-011,
  6.040734e-014, 1.360983e-015, 1.872597e-012, -3.143038e-012,
  1.797076e-013, -9.079147e-015, -1.076987e-012, 3.060381e-011,
  6.825358e-014, -2.041189e-015, 2.365594e-012, -4.178561e-012,
  1.182966e-013, -1.460926e-015, 6.089823e-013, 3.217946e-011,
  7.627887e-014, -1.547783e-015, 2.728722e-013, -6.050241e-012,
  1.200153e-013, -3.894285e-015, 2.681911e-013, 3.09202e-011,
  7.713833e-014, -4.13596e-015, 1.998096e-014, -6.617119e-012,
  1.292035e-013, -5.463726e-015, 1.46528e-012, 3.236806e-011,
  7.855043e-014, -7.587312e-015, -5.314556e-013, -9.95334e-012,
  1.372709e-013, -7.731402e-015, 1.099422e-012, 3.404178e-011,
  8.45996e-014, -1.662075e-015, -2.645254e-014, -9.575007e-012,
  1.401064e-013, -6.730165e-015, -1.244318e-012, 3.272412e-011,
  8.737055e-014, -3.46151e-015, -4.026754e-013, -8.021222e-012,
  1.428225e-013, -7.080293e-015, 1.487418e-012, 3.426416e-011,
  9.293358e-014, -6.350124e-015, -1.097792e-012, -1.089647e-011,
  1.527196e-013, -6.898272e-015, 1.155808e-012, 3.84202e-011,
  -2.114002e-014, 1.244478e-014, 2.026458e-012, -5.812541e-012,
  2.306213e-013, -1.860104e-014, 1.385241e-012, 4.090168e-011,
  1.019832e-013, -5.215632e-015, 3.364835e-012, -3.921263e-012,
  1.669549e-013, -7.970613e-015, -2.515199e-013, 4.03697e-011,
  1.012803e-013, -5.124378e-015, -9.25557e-012, -2.065976e-011,
  1.737355e-013, -1.253589e-014, 1.64842e-012, 4.321789e-011,
  1.134815e-013, 1.540177e-015, -5.818735e-012, -1.464718e-011,
  1.826885e-013, -1.081203e-014, 1.961012e-011, 5.55872e-011,
  1.047993e-013, 8.843506e-017, 9.605036e-012, 2.155091e-012,
  2.555773e-013, -1.860648e-014, 4.519798e-012, 5.278734e-011,
  1.236854e-013, -4.985132e-015, 2.817799e-012, -8.829189e-012,
  2.1714e-013, -1.300632e-014, 7.738336e-012, 5.364023e-011,
  1.345503e-013, -1.503284e-015, -2.533084e-012, -1.42537e-011,
  2.169246e-013, -5.404516e-015, -7.81961e-012, 4.826787e-011,
  1.381239e-013, -4.798667e-016, -1.427027e-013, -1.16602e-011,
  2.202342e-013, -8.287701e-015, 2.639632e-014, 5.348944e-011,
  1.009364e-013, 2.490405e-015, -3.103602e-012, -1.495735e-011,
  2.196856e-013, -5.039661e-015, 2.40119e-012, 5.9967e-011,
  8.924084e-014, 6.831865e-015, -1.765583e-012, -1.372674e-011,
  2.480853e-013, -8.606077e-015, 5.820068e-012, 6.418653e-011,
  1.602338e-013, -4.067726e-015, 7.756363e-013, -1.490969e-011,
  2.647708e-013, -2.22537e-015, 3.222396e-012, 6.966117e-011,
  1.75105e-013, -2.116636e-015, -2.157006e-013, -1.710295e-011,
  2.8004e-013, 4.99215e-015, -1.308971e-012, 7.157551e-011,
  1.706274e-013, 4.205388e-016, 1.125956e-012, -1.644553e-011,
  2.979836e-013, -2.64968e-015, 8.676566e-012, 7.798252e-011,
  1.782367e-013, -7.970932e-015, -8.914109e-012, -2.515257e-011,
  3.155262e-013, -1.62496e-014, 1.090842e-011, 8.186497e-011,
  2.019608e-013, -1.152222e-014, -2.154044e-012, -1.958846e-011,
  3.414201e-013, -2.449983e-014, -1.856826e-012, 8.349867e-011,
  2.087699e-013, -1.483075e-014, -2.901376e-012, -2.003154e-011,
  3.48174e-013, -1.230862e-014, 1.227766e-011, 9.754331e-011,
  2.202486e-013, -3.591038e-015, -5.465183e-012, -2.449647e-011,
  3.717067e-013, -2.316929e-015, 1.204963e-011, 1.00798e-010,
  1.315322e-013, 1.026687e-014, 1.074401e-012, -2.110691e-011,
  2.816286e-013, 1.398014e-014, 1.031258e-011, 1.107593e-010,
  2.474265e-013, 1.046868e-015, 8.29181e-012, -1.248353e-011,
  4.216813e-013, -9.347885e-015, 1.027818e-011, 1.11134e-010,
  2.628918e-013, -8.455748e-015, 6.937916e-013, -2.847115e-011,
  4.61662e-013, -1.120409e-014, 1.849702e-011, 1.306016e-010,
  2.807375e-013, -7.068625e-015, -7.476161e-012, -3.149235e-011,
  4.879192e-013, -2.182075e-014, 6.796342e-012, 1.23915e-010,
  2.226041e-013, 4.889158e-015, -8.832453e-012, -3.472515e-011,
  5.293425e-013, -1.89297e-014, 3.265815e-012, 1.305353e-010,
  3.177356e-013, -1.282719e-014, -8.737794e-012, -3.813694e-011,
  5.674857e-013, -2.151257e-014, 6.390754e-012, 1.403636e-010,
  3.527044e-013, -1.87729e-014, -9.876722e-012, -4.257108e-011,
  6.098346e-013, -3.170482e-014, 6.857832e-012, 1.481733e-010,
  3.844124e-013, -3.397178e-014, -1.429074e-011, -5.900141e-011,
  6.564463e-013, -4.346943e-014, 1.506646e-011, 1.73195e-010,
  4.172338e-013, -2.519673e-014, 5.418664e-012, -2.881212e-011,
  7.706528e-013, -4.041317e-014, 2.39596e-011, 1.887532e-010,
  4.576898e-013, -2.397996e-014, -3.717464e-012, -5.222697e-011,
  8.081822e-013, -4.261153e-014, 1.453319e-011, 1.813957e-010,
  4.895959e-013, -1.825668e-014, 4.592466e-012, -5.077009e-011,
  8.32896e-013, -1.336621e-014, 2.422924e-011, 2.108748e-010,
  5.459229e-013, -9.472764e-015, -1.344443e-011, -6.846332e-011,
  9.145983e-013, -2.083938e-014, -2.561251e-013, 2.050109e-010,
  5.964282e-013, -1.236606e-014, 9.169158e-012, -5.172202e-011,
  9.966102e-013, -1.399271e-014, 4.397186e-012, 2.180544e-010,
  6.582538e-013, -1.829346e-014, -9.157442e-012, -8.704881e-011,
  1.076327e-012, -4.144125e-014, 9.261336e-012, 2.456322e-010,
  7.307679e-013, -1.916381e-014, -4.964579e-012, -9.840757e-011,
  1.164561e-012, -3.727298e-014, 1.306165e-011, 2.758163e-010,
  8.160262e-013, -1.746131e-014, -2.038512e-012, -1.143995e-010,
  1.257979e-012, -2.342775e-014, 6.64117e-012, 3.066763e-010,
  9.050707e-013, -1.61385e-014, -4.990532e-012, -1.377458e-010,
  1.358241e-012, -2.078428e-014, 5.718666e-012, 3.474219e-010,
  1.013104e-012, -1.618746e-014, 2.725378e-012, -1.533074e-010,
  1.465185e-012, -2.12565e-014, 3.090323e-012, 3.914999e-010,
  1.129768e-012, 2.385275e-016, -1.169656e-013, -1.79144e-010,
  1.566411e-012, -3.749735e-015, -3.0949e-013, 4.534408e-010,
  1.238424e-012, 1.371574e-014, 2.510452e-012, -2.026294e-010,
  1.676103e-012, 1.727468e-014, -3.076559e-012, 5.26833e-010,
  1.421823e-012, -3.266454e-015, -1.292309e-011, -2.588414e-010,
  1.720567e-012, 3.675195e-014, -2.641147e-011, 5.723043e-010,
  1.507166e-012, -6.195256e-015, 4.709614e-011, -2.416208e-010,
  1.891009e-012, 1.7821e-014, 1.29785e-010, 7.978286e-010,
  1.587579e-012, 5.217959e-016, 2.770977e-011, -2.067488e-010,
  2.058676e-012, 1.989217e-015, 1.898432e-011, 8.868271e-010,
  1.69658e-012, -1.761091e-015, 2.462238e-011, -1.849721e-010,
  2.252065e-012, -1.546586e-014, 1.116985e-012, 1.054766e-009,
  1.704711e-012, -7.539542e-015, -4.102209e-013, -1.947165e-010,
  2.379051e-012, 7.221262e-015, 9.999273e-012, 1.25582e-009,
  1.67308e-012, -2.350824e-014, 2.809624e-012, -1.136247e-010,
  2.606305e-012, -3.180108e-014, 2.631534e-011, 1.498851e-009,
  1.544481e-012, -7.028866e-014, -2.093005e-012, 2.593755e-011,
  2.929531e-012, -9.142559e-014, 5.377721e-011, 1.771915e-009,
  1.275126e-012, -4.955752e-014, 4.496696e-012, 2.332511e-010,
  3.387296e-012, -9.020855e-014, 4.849566e-011, 2.071187e-009,
  8.187526e-013, -3.140906e-014, 6.870359e-012, 5.488426e-010,
  4.07239e-012, -1.040459e-013, 5.553185e-011, 2.402914e-009,
  1.833316e-013, -1.918879e-014, 1.043601e-011, 1.003726e-009,
  5.132555e-012, -1.725662e-013, 7.550355e-011, 2.731662e-009,
  -7.658714e-013, -1.356219e-014, 1.999652e-011, 1.63352e-009,
  6.759477e-012, -3.247616e-013, 1.119039e-010, 3.026495e-009,
  -2.014898e-012, -2.602584e-015, 4.507892e-011, 2.490693e-009,
  9.241378e-012, -5.255626e-013, 1.497057e-010, 3.231138e-009,
  -3.646568e-012, 1.227432e-014, 6.848506e-011, 3.60034e-009,
  1.299218e-011, -8.482273e-013, 1.994903e-010, 3.26696e-009,
  -5.600457e-012, 1.402061e-014, 1.117431e-010, 5.023111e-009,
  1.870405e-011, -1.262387e-012, 2.097853e-010, 2.961727e-009,
  -7.527454e-012, -6.211988e-014, 1.798359e-010, 6.773735e-009,
  2.727699e-011, -2.203276e-012, 2.857348e-010, 2.210025e-009,
  -9.016726e-012, -3.284875e-013, 2.764507e-010, 8.840586e-009,
  3.999469e-011, -3.544193e-012, 3.483652e-010, 6.708916e-010,
  -8.04482e-012, -8.510963e-013, 3.299576e-010, 1.118977e-008,
  5.875379e-011, -4.699583e-012, 3.077341e-010, -2.007533e-009,
  -4.763413e-012, -2.003606e-012, 3.879328e-010, 1.358815e-008,
  8.755643e-011, -6.726461e-012, 2.586479e-010, -6.483517e-009,
  6.881907e-012, -4.56371e-012, 4.800257e-010, 1.555446e-008,
  1.2984e-010, -1.02511e-011, 2.592836e-010, -1.375332e-008,
  3.227664e-011, -8.100827e-012, 4.951973e-010, 1.60908e-008,
  1.938308e-010, -1.351624e-011, 1.937647e-010, -2.517955e-008,
  8.773585e-011, -1.373015e-011, 4.001383e-010, 1.314451e-008,
  2.884234e-010, -1.653098e-011, 1.224751e-010, -4.259132e-008,
  2.030932e-010, -2.187194e-011, 2.367023e-010, 2.460427e-009,
  4.355033e-010, -1.900889e-011, 1.795434e-010, -6.976097e-008,
  4.427074e-010, -3.435313e-011, 1.586847e-010, -2.490446e-008,
  6.629829e-010, -1.921556e-011, 7.362406e-010, -1.115506e-007,
  9.51325e-010, -6.687108e-011, 1.021553e-009, -9.141423e-008,
  1.015279e-009, -1.995666e-011, 3.107314e-009, -1.780041e-007,
  1.961923e-009, -1.382554e-010, 5.693817e-009, -2.564169e-007,
  1.537139e-009, -1.877268e-011, 8.500514e-009, -2.870447e-007,
  2.906412e-009, -3.209273e-010, 2.477005e-008, -7.023682e-007,
  2.044687e-009, -1.175972e-011, 2.015833e-008, -4.741695e-007,
  -2.4371e-009, -6.530367e-010, 8.588849e-008, -1.824169e-006,
  1.708062e-009, 3.948053e-013, 4.099665e-008, -7.693349e-007,
  -1.241482e-008, -6.907303e-010, 1.443044e-007, -3.176909e-006,
  1.55214e-009, 3.249477e-011, 5.120048e-008, -1.012575e-006,
  -1.446957e-008, -6.646975e-010, 1.473276e-007, -3.579323e-006,
  1.636457e-009, 1.509586e-012, 4.388047e-008, -1.067093e-006,
  -1.142095e-008, -1.058721e-009, 9.884732e-008, -2.983462e-006,
  2.015712e-009, -1.103432e-010, 2.834157e-008, -9.054936e-007,
  -1.019035e-009, -1.128542e-009, 3.714581e-008, -1.614246e-006,
  2.546288e-009, -1.0595e-010, 1.587618e-008, -6.137018e-007,
  3.019229e-009, -4.620312e-010, 1.018115e-008, -6.153744e-007,
  1.997231e-009, -4.023641e-011, 8.699915e-009, -3.950069e-007,
  1.867956e-009, -1.046874e-010, 2.488968e-009, -2.294153e-007,
  1.384845e-009, -7.032847e-012, 3.496032e-009, -2.523402e-007,
  9.036636e-010, -1.961647e-011, 3.189959e-010, -8.400105e-008,
  9.201224e-010, -3.62841e-012, 9.751403e-010, -1.614474e-007,
  4.275895e-010, -1.54172e-011, 1.138217e-010, -2.368089e-008,
  6.071609e-010, -1.084054e-011, 2.567876e-010, -1.031007e-007,
  2.005476e-010, -1.550066e-011, 1.05494e-010, 1.522156e-009,
  4.056461e-010, -1.730197e-011, 7.539842e-011, -6.562602e-008,
  9.069033e-011, -1.474134e-011, 3.538689e-010, 1.152812e-008,
  2.743014e-010, -2.04023e-011, 1.457684e-010, -4.140927e-008,
  3.615639e-011, -1.01834e-011, 6.679923e-010, 1.494257e-008,
  1.862356e-010, -1.60167e-011, 4.119178e-010, -2.516306e-008,
  9.605995e-012, -5.211043e-012, 4.048578e-010, 1.454771e-008,
  1.272622e-010, -1.016149e-011, 5.005522e-010, -1.450349e-008,
  -2.162775e-012, -2.071152e-012, 2.507618e-010, 1.30869e-008,
  8.747972e-011, -5.157054e-012, 4.299601e-010, -7.584714e-009,
  -7.040785e-012, -1.075169e-012, 1.857139e-010, 1.099644e-008,
  6.009613e-011, -3.994755e-012, 5.102611e-010, -3.030875e-009,
  -8.714827e-012, -5.78406e-013, 1.357148e-010, 8.918349e-009,
  4.171963e-011, -2.872813e-012, 4.80725e-010, -2.882026e-010,
  -7.810396e-012, -3.512025e-013, 1.057922e-010, 7.026517e-009,
  2.898154e-011, -2.319121e-012, 4.433787e-010, 1.330781e-009,
  -6.24319e-012, -2.848564e-013, -2.188178e-011, 5.257444e-009,
  2.023094e-011, -1.619086e-012, 3.705649e-010, 2.274285e-009,
  -4.604588e-012, -2.111136e-013, -9.785323e-012, 4.01453e-009,
  1.425892e-011, -7.182915e-013, 2.15553e-010, 2.700881e-009,
  -3.034993e-012, -1.634594e-013, -5.27082e-011, 2.911583e-009,
  1.018916e-011, -2.989316e-014, 7.041402e-011, 2.838658e-009,
  -1.707752e-012, -1.212912e-013, -7.202325e-011, 2.004397e-009,
  7.432485e-012, -4.397328e-014, 2.810536e-011, 2.722596e-009,
  -6.84799e-013, -1.392386e-013, -2.055992e-011, 1.36428e-009,
  5.577841e-012, -1.394725e-013, 6.946783e-011, 2.560778e-009,
  2.185818e-014, -3.134238e-013, -2.499473e-010, 5.047794e-010,
  4.28317e-012, -3.08983e-013, 1.195169e-010, 2.462367e-009,
  5.8339e-013, -2.705925e-013, -4.63743e-010, -2.076284e-010,
  3.433166e-012, -5.246189e-013, 7.069985e-011, 2.173062e-009,
  9.55905e-013, -1.470684e-013, 1.069797e-011, 2.19641e-010,
  2.934378e-012, 1.018305e-015, -1.286644e-010, 1.524232e-009,
  1.179177e-012, 6.602385e-014, -1.272066e-010, -1.429035e-010,
  2.448893e-012, -1.925367e-013, -1.198715e-010, 1.33847e-009,
  1.319645e-012, 2.65221e-014, 3.418427e-012, -6.877775e-011,
  2.267519e-012, -3.755714e-014, -2.851568e-011, 1.261717e-009,
  1.375662e-012, 2.643323e-014, 6.133048e-011, -4.04278e-011,
  2.092725e-012, 5.447487e-014, -3.122885e-011, 1.078633e-009,
  1.357564e-012, -6.370126e-014, -1.166068e-011, -1.988291e-010,
  1.92621e-012, -7.479295e-015, 4.443229e-011, 1.049761e-009,
  1.304005e-012, -1.126445e-013, 2.264997e-011, -1.499202e-010,
  1.798591e-012, 6.140647e-014, 1.132123e-010, 1.002603e-009,
  1.253574e-012, 3.903218e-014, 1.01766e-010, -4.057344e-011,
  1.699804e-012, 9.82344e-014, -1.773225e-011, 6.540217e-010,
  1.173284e-012, -2.509024e-015, 1.178414e-011, -1.809539e-010,
  1.578035e-012, -1.192923e-014, -4.893841e-012, 5.887814e-010,
  1.083538e-012, -1.927157e-014, 2.872463e-012, -1.845203e-010,
  1.484554e-012, -2.774347e-014, 1.586572e-011, 5.211627e-010,
  9.932067e-013, -2.04904e-014, -3.218417e-011, -2.218783e-010,
  1.38631e-012, -2.506422e-014, 1.801569e-011, 4.67058e-010,
  9.116948e-013, 5.797803e-015, 6.18317e-012, -1.48554e-010,
  1.303233e-012, 3.303461e-014, -2.721823e-013, 3.967395e-010,
  8.211091e-013, 2.626725e-014, 1.617517e-011, -1.201391e-010,
  1.220499e-012, 5.054904e-014, -2.597043e-012, 3.432701e-010,
  7.452329e-013, 3.197598e-014, 2.441068e-011, -9.75709e-011,
  1.14364e-012, 5.458995e-014, -2.262484e-011, 2.741962e-010,
  6.997734e-013, 2.77728e-014, 5.125947e-011, -3.517329e-011,
  1.043243e-012, 3.652356e-014, -1.642868e-011, 2.494165e-010,
  6.095797e-013, -3.383881e-014, 1.797167e-011, -5.733349e-011,
  9.892047e-013, 4.13377e-015, 4.230232e-011, 3.00158e-010,
  5.620634e-013, -1.223754e-014, -6.693674e-011, -2.165866e-010,
  9.017343e-013, -1.48702e-013, -5.468561e-011, 1.277287e-010,
  4.759504e-013, -1.802047e-013, -1.429238e-010, -3.013131e-010,
  8.292867e-013, -1.897415e-013, 8.132059e-011, 3.472714e-010,
  4.628269e-013, 5.102386e-014, -1.675622e-010, -3.683277e-010,
  7.011558e-013, -6.00719e-013, -1.995565e-010, -1.222748e-010,
  5.789488e-013, 1.614933e-013, 6.179429e-012, -8.274209e-011,
  7.202973e-013, -2.004659e-014, -1.786602e-010, -1.234943e-010,
  3.704723e-013, -4.947032e-014, -1.304362e-010, -2.115586e-010,
  6.205195e-013, -3.72719e-013, 1.396237e-010, 3.83156e-010,
  3.774553e-013, 1.495283e-013, -3.979403e-010, -7.502367e-010,
  5.480104e-013, -5.850427e-013, -1.483576e-010, -5.655363e-011,
  3.230442e-013, 1.720548e-014, -8.025166e-011, -1.801247e-010,
  5.854028e-013, -8.733852e-014, -2.012363e-011, 9.282924e-011,
  3.468597e-013, 1.983394e-014, -5.214329e-011, -1.499143e-010,
  4.785519e-013, -5.586294e-014, -3.589324e-011, 6.537828e-011,
  2.880239e-013, -1.014767e-015, -2.658079e-011, -8.679266e-011,
  4.978156e-013, -5.578773e-014, -9.065733e-012, 8.436404e-011,
  2.635603e-013, -1.339395e-014, 2.448412e-011, 3.139527e-011,
  4.868487e-013, -4.090157e-015, -2.320449e-013, 1.042661e-010,
  2.374757e-013, -5.087663e-014, -6.343844e-012, -1.247255e-011,
  4.494263e-013, -4.861972e-014, 5.2922e-011, 1.895224e-010,
  1.808361e-013, -8.771312e-014, -1.226905e-010, -2.179545e-010,
  3.655097e-013, -1.691368e-013, 1.910046e-011, 1.240216e-010,
  1.85714e-013, -4.924105e-014, 5.645924e-012, 1.50754e-012,
  3.87589e-013, -3.253058e-014, 9.653885e-012, 1.2022e-010,
  1.996569e-013, -1.093868e-013, 1.285364e-010, 2.127286e-010,
  3.984568e-013, 1.246522e-013, 1.249583e-010, 2.484002e-010,
  2.0017e-013, 2.378074e-015, 4.127627e-011, 5.205622e-011,
  3.524885e-013, -7.698821e-015, -9.984678e-012, 5.155127e-011,
  1.755814e-013, -5.917821e-014, 1.304538e-010, 1.648894e-010,
  3.258713e-013, 2.066622e-014, -3.32913e-011, 1.499346e-012,
  1.374496e-013, -9.87938e-014, 9.636657e-011, 1.507578e-010,
  3.284753e-013, 6.283923e-014, 1.146596e-010, 2.391391e-010,
  1.849301e-013, 1.776245e-013, 4.784264e-010, 7.267968e-010,
  3.389649e-013, 2.047515e-013, -1.061738e-010, -1.43954e-010,
  1.80254e-013, 1.354133e-013, -2.91187e-011, -8.200753e-011,
  2.772578e-013, -3.366747e-014, -1.637165e-010, -1.652923e-010,
  8.815209e-014, -3.940461e-013, 1.70939e-010, 2.848539e-010,
  3.358042e-013, 3.492043e-013, 2.775311e-010, 5.445463e-010,
  1.364129e-013, -3.288518e-013, -1.141946e-010, -1.834464e-010,
  3.798972e-013, -1.120274e-013, 2.738845e-010, 5.317827e-010,
  1.658029e-013, 1.42112e-013, 2.137318e-010, 3.020517e-010,
  2.580781e-013, 1.365998e-013, -9.057295e-011, -1.201399e-010,
  1.026798e-013, -2.169014e-013, -1.231273e-010, -1.718256e-010,
  2.001521e-013, -1.339758e-013, 1.756823e-010, 3.541484e-010,
  1.404315e-013, 8.134929e-014, 5.60321e-010, 9.031542e-010,
  2.919845e-013, 4.552712e-013, 4.737761e-011, 2.278719e-011,
  1.90414e-013, -5.849668e-014, 1.266758e-012, 4.758628e-012,
  2.42173e-013, -4.583886e-014, -1.340549e-012, 3.374652e-011,
  1.086198e-013, -5.669483e-014, -1.529003e-011, -1.409038e-011,
  2.013221e-013, -6.301218e-014, 4.481032e-011, 9.42857e-011,
  6.49355e-014, -2.369065e-013, -3.295011e-011, -2.58753e-011,
  1.795583e-013, -3.813694e-014, 2.077578e-010, 3.701686e-010,
  8.207776e-014, -1.28385e-013, 5.473989e-011, 1.084482e-010,
  1.916404e-013, 4.940762e-014, 1.251372e-010, 2.263667e-010,
  1.34126e-013, -9.51997e-015, 2.91132e-011, 4.254733e-011,
  1.204049e-013, -8.230329e-015, -4.008414e-012, 2.457809e-011,
  1.015075e-013, -1.831064e-014, 1.448618e-012, -1.147299e-011,
  1.403681e-013, -3.09723e-014, -2.945459e-012, 2.976297e-011,
  8.594805e-014, -1.74285e-014, 4.58261e-012, -7.469939e-012,
  1.549353e-013, -2.121057e-014, 1.324532e-011, 4.907449e-011,
  8.206666e-014, -1.958995e-014, -6.096598e-012, -2.162011e-011,
  1.462341e-013, -3.03548e-014, 1.179199e-011, 3.553826e-011,
  7.528919e-014, -4.280593e-014, -8.186091e-011, -1.508903e-010,
  1.302996e-013, -1.054067e-013, -6.790172e-012, 4.257176e-011,
  6.822298e-014, -9.675014e-014, 2.332506e-011, 4.879667e-011,
  1.416648e-013, 9.412902e-015, 9.490457e-011, 1.800068e-010,
  8.548908e-014, 6.417759e-014, -2.549475e-011, -6.149248e-011,
  1.200021e-013, -7.282934e-014, -5.429661e-011, -7.79484e-011,
  6.508327e-014, -6.432389e-014, 1.536103e-011, 1.954766e-011,
  1.267699e-013, -2.005714e-015, 5.189824e-011, 1.136038e-010,
  6.108703e-014, 1.013287e-013, 3.270646e-011, 3.824163e-011,
  1.264196e-013, 1.5037e-014, -5.407164e-011, -7.027106e-011,
  -4.523934e-014, 9.655882e-014, -6.146023e-011, -1.452906e-010,
  1.686607e-013, -1.090462e-013, -6.493722e-012, 4.688492e-011,
  2.504613e-014, -2.325284e-013, -2.433447e-010, -3.988138e-010,
  8.32527e-014, -2.076924e-013, 1.7837e-010, 3.52324e-010,
  1.022556e-013, -5.65766e-014, -1.123243e-010, -1.463093e-010,
  1.188759e-013, 8.737532e-014, 7.831732e-011, 1.99989e-010,
  1.381002e-013, -2.436608e-013, 3.324072e-010, 6.669479e-010,
  4.711092e-014, 4.854997e-013, 4.758072e-010, 8.205319e-010,
  1.041621e-013, 3.532666e-013, -1.928917e-010, -3.32809e-010,
  7.778131e-014, -5.692101e-013, -3.841973e-010, -6.740459e-010,
  2.335466e-014, 9.939806e-014, -3.651374e-010, -5.96187e-010,
  1.412292e-014, -6.866287e-013, -1.721116e-010, -2.837316e-010,
  3.197427e-013, 3.731871e-013, 2.769569e-010, 4.939198e-010,
  -5.576236e-014, -8.430069e-013, 2.813736e-010, 5.093367e-010,
  1.502957e-013, 9.221923e-015, 4.318803e-013, 4.643146e-011,
  1.109707e-014, 2.359742e-014, 6.803675e-011, 1.836709e-010,
  1.807198e-013, -4.119261e-013, 2.939585e-010, 4.881806e-010,
  2.773731e-013, 4.208169e-013, 5.177019e-010, 8.907657e-010,
  -9.280666e-015, 1.051478e-014, 1.262134e-010, 1.945358e-010,
  1.904779e-013, 1.637743e-013, -1.60447e-011, -9.1208e-011,
  2.510131e-013, -8.319791e-014, 6.980827e-011, 3.57316e-010,
  -2.198685e-013, -5.517298e-015, 1.578764e-010, 4.177413e-010,
  -2.153575e-013, -6.583055e-014, -2.146772e-011, -1.630993e-010,
  3.048574e-013, 2.172446e-014, -5.016041e-011, -2.227395e-010,
  -4.116965e-013, -1.862271e-013, -1.169471e-010, -5.40841e-010,
  1.023274e-012, 2.388687e-013, 9.633741e-011, -9.307063e-011,
  -1.569817e-013, 5.965707e-014, -8.660261e-011, -3.392941e-010,
  4.290389e-013, -9.640223e-014, -2.189829e-010, -4.415556e-010,
  1.695984e-013, -1.840317e-013, -2.485425e-010, -5.306772e-010,
  3.049446e-013, -1.406142e-013, 7.999893e-011, 2.264927e-010,
  -3.306831e-013, 9.607346e-014, -3.551326e-010, -7.39591e-010,
  1.597656e-013, -3.567088e-013, -5.134735e-010, -9.809352e-010,
  -6.616355e-015, -1.751062e-014, 7.332231e-011, 1.096692e-010,
  6.818673e-014, 9.651816e-015, -2.399111e-011, -5.253378e-011,
  6.627538e-014, -8.354232e-014, -3.065026e-011, -1.387462e-010,
  2.533848e-013, 3.381547e-014, 9.118813e-011, 1.828653e-010,
  -3.843049e-013, 8.475923e-014, 3.754319e-010, 8.233375e-010,
  -2.629543e-013, 1.454711e-013, -1.595098e-010, -4.788083e-010,
  8.941527e-015, -1.110571e-014, 4.12552e-011, 5.785167e-011,
  4.949256e-014, -5.602527e-015, 1.730522e-011, 1.563679e-011,
  2.312873e-014, -2.483268e-014, -4.380222e-011, -6.235273e-011,
  4.422033e-014, -5.548641e-014, 2.53304e-011, 5.685964e-011,
  -1.045594e-013, -9.523581e-015, -6.996641e-011, -1.693836e-010,
  1.399983e-013, -6.243059e-014, -4.072315e-011, -8.296739e-011,
  2.630401e-014, -6.490524e-014, -5.519419e-011, -1.016626e-010,
  4.45945e-014, -4.988676e-014, 5.373019e-011, 1.09728e-010,
  2.903224e-014, -4.783539e-015, -9.683068e-012, -2.330484e-011,
  5.855895e-014, -1.876607e-014, -1.898462e-013, 5.732144e-012,
  2.516474e-014, -6.67902e-015, 2.696641e-012, -4.850118e-012,
  4.93808e-014, -1.912375e-014, -3.894711e-012, -7.956e-012,
  2.333846e-014, -1.254391e-014, 3.866858e-012, -5.63825e-013,
  4.426398e-014, -1.83841e-014, 7.070344e-012, 1.371866e-011,
  2.253526e-014, -7.558593e-015, 4.113792e-012, -2.74523e-012,
  4.568033e-014, -3.445718e-014, 1.766808e-012, 9.70944e-012,
  2.584745e-014, -9.814521e-015, -3.188057e-013, -8.74935e-013,
  4.416877e-014, -2.197281e-014, 1.499463e-012, 6.284145e-012,
  2.395317e-014, -9.996857e-015, 1.247521e-012, -1.001229e-011,
  2.660262e-014, -3.248088e-014, 4.735592e-012, 5.43589e-012,
  -3.587329e-014, -9.997665e-015, -2.565127e-011, -4.063128e-011,
  1.712407e-014, -4.256825e-014, 7.710187e-013, 1.436713e-011,
  -7.396932e-015, 1.15824e-014, 4.942514e-011, 8.998786e-011,
  5.325154e-014, 3.592417e-014, -5.204961e-012, -1.291097e-011,
  5.309332e-014, 1.231968e-013, 7.301659e-011, 1.051717e-010,
  5.541558e-014, 4.227199e-014, -1.024906e-010, -1.857734e-010,
  2.232873e-014, -4.656037e-014, -9.812591e-012, -1.922766e-011,
  3.447196e-014, -1.813123e-014, 4.712377e-011, 9.876944e-011,
  -4.529213e-015, -2.468565e-014, 1.448103e-011, 2.181121e-011,
  6.352303e-014, -1.083457e-014, 1.650321e-011, 4.275464e-011,
  -4.135445e-014, -2.729284e-014, 5.457925e-011, 1.143555e-010,
  2.702357e-014, -2.180965e-014, -6.853043e-012, -6.262573e-012,
  6.447235e-014, -1.404318e-014, 2.093873e-011, 8.276413e-011,
  -3.226564e-014, 1.956348e-015, 3.785466e-011, 8.459597e-011,
  -3.40115e-014, -2.624603e-015, -4.472639e-011, -9.19525e-011,
  1.032308e-013, -2.191693e-014, -5.182122e-011, -1.192388e-010,
  1.773439e-013, -2.387418e-014, -1.156031e-010, -2.205526e-010,
  1.117544e-013, -3.310721e-014, 9.524141e-011, 2.680846e-010,
  -7.916237e-013, 7.665654e-014, -6.320458e-011, -2.454102e-010,
  3.085709e-013, 4.140715e-014, -4.086797e-010, -1.010589e-009,
  1.751315e-013, -3.363067e-014, 5.626567e-011, 1.384615e-010,
  -7.67534e-014, 1.070064e-014, 1.489273e-010, 3.498392e-010,
  -1.951723e-014, -7.493852e-015, 1.559919e-010, 3.490571e-010,
  -1.415843e-013, 1.983657e-014, -1.278659e-011, -6.872437e-011,
  -7.180386e-015, -1.045593e-014, -3.00123e-011, -1.204872e-010,
  7.220444e-014, 4.458295e-015, 6.689482e-011, 9.498128e-011,
  -4.144585e-013, 7.039229e-014, -3.868024e-010, -1.016721e-009,
  8.255455e-013, -1.217528e-013, -2.17825e-010, -5.252058e-010,
  -6.006871e-014, 5.988606e-014, -1.80294e-010, -4.781072e-010,
  3.697028e-013, -3.576728e-014, -1.774908e-010, -3.454621e-010,
  -1.343252e-013, 7.805454e-015, 1.805612e-010, 3.212636e-010,
  -1.672698e-014, 8.815569e-014, -9.342845e-011, -2.258956e-010,
  1.125692e-013, 1.485782e-014, -9.886631e-011, -2.985233e-010,
  1.757235e-013, -2.435052e-014, -2.088722e-011, 7.661662e-011,
  -3.538601e-013, 1.459183e-013, -4.289051e-010, -1.1458e-009,
  6.88737e-013, -3.291389e-014, -4.152312e-010, -9.315353e-010,
  3.061581e-013, 1.384246e-013, -4.489409e-011, -1.434566e-010,
  1.771331e-013, 2.858843e-014, 1.684966e-010, 5.255379e-010,
  8.479666e-013, -2.241051e-013, 1.624256e-011, 3.174505e-011,
  1.792748e-014, 7.45439e-014, 6.847471e-010, 1.741738e-009,
  -4.087179e-013, -2.741123e-013, -9.364387e-010, -1.837873e-009,
  3.537162e-013, -6.1587e-013, -1.166749e-010, -2.823601e-010,
  -4.612037e-013, 6.440346e-013, -1.628614e-010, -2.670959e-010,
  -2.763088e-013, -3.774577e-013, -8.552963e-010, -1.506905e-009,
  6.554374e-014, 8.64883e-014, -1.172165e-010, -2.605851e-010,
  9.996554e-014, -1.216942e-013, -1.462831e-010, -2.46704e-010,
  1.402534e-013, -3.033738e-014, -6.273933e-011, -1.291631e-010,
  -3.331957e-014, -1.070413e-013, 6.594254e-011, 2.10427e-010,
  3.232407e-014, 1.872299e-014, -3.190497e-011, -2.384378e-011,
  -7.488254e-014, -4.799258e-014, 8.006614e-012, 1.240685e-011,
  1.572645e-013, -2.350107e-014, 1.224583e-011, 8.312189e-011,
  -7.037317e-014, 1.380168e-014, 1.081349e-010, 2.67317e-010,
  6.913806e-014, -1.91712e-014, -2.682611e-011, -3.045147e-011,
  -6.443428e-014, -3.907716e-015, 3.034532e-011, 8.450911e-011,
  -1.009685e-014, -1.046334e-014, -1.354109e-011, 1.001359e-011,
  -6.527719e-015, -7.494554e-015, -9.992618e-012, -1.321989e-011,
  -1.301988e-014, -1.002462e-014, 2.733352e-011, 2.976839e-011,
  3.595569e-014, -1.533734e-014, 2.763214e-013, -9.556291e-012,
  -1.066335e-014, -1.678751e-014, 1.426667e-011, 2.338364e-011,
  1.759538e-014, -2.356418e-014, 1.793963e-011, 1.358287e-011,
  -6.216594e-014, 7.02783e-015, 1.453718e-011, 2.180095e-011,
  -2.227026e-014, -9.706385e-015, 1.110388e-011, 1.007867e-011,
  1.901953e-014, -5.059241e-015, -7.733532e-013, -1.677276e-011,
  1.527137e-014, -2.109787e-014, 2.823683e-011, 3.450215e-011,
  1.533736e-013, -2.604441e-014, -7.602175e-011, -1.72753e-010,
  9.92344e-014, -1.013694e-013, 1.212933e-010, 2.739203e-010,
  8.393844e-014, -5.464016e-014, 1.674554e-010, 2.449687e-010,
  7.524138e-014, -1.090948e-013, 1.386754e-010, 3.316481e-010,
  -6.901249e-015, 9.547103e-014, -6.64919e-011, -1.024446e-010,
  -1.621554e-014, -1.05054e-013, -2.072759e-010, -3.609493e-010,
  1.026897e-013, 2.609075e-013, 2.987343e-011, 6.014131e-011,
  -4.764086e-014, -1.087173e-014, -2.058339e-010, -3.439714e-010,
  9.939067e-014, 1.514976e-013, 4.929748e-011, 9.771246e-011,
  -8.760661e-014, -6.408233e-015, -1.59224e-010, -2.537044e-010,
  -2.494963e-013, -1.642085e-013, 1.549399e-010, 5.676571e-010,
  -2.802483e-013, 1.388077e-013, -9.902686e-011, -2.762049e-010,
  -7.483553e-013, 6.756965e-015, -1.204938e-010, -3.185888e-010,
  3.154208e-013, -5.020179e-014, -4.194685e-010, -1.172924e-009,
  -1.23838e-013, -6.555829e-015, -3.601186e-010, -8.408e-010,
  4.725528e-013, -1.83748e-013, -3.913529e-012, -1.342689e-010,
  6.015442e-014, -9.337861e-014, -2.129512e-010, -5.18719e-010,
  3.462257e-013, -3.060096e-014, 1.476713e-010, 2.439179e-010,
  1.088628e-013, 1.490235e-013, 4.604571e-011, 9.567377e-011,
  -1.843213e-014, -4.106367e-014, -1.783539e-010, -2.605897e-010,
  1.245235e-013, -2.154127e-014, 1.030551e-010, 2.498076e-010,
  -1.878543e-013, -3.360536e-014, -1.137253e-011, 8.58843e-012,
  6.779305e-013, -5.883856e-014, 2.064066e-010, 4.376794e-010,
  -2.211711e-013, -9.898571e-015, 3.417387e-010, 8.742359e-010,
  3.310879e-015, 4.932279e-014, 3.559043e-010, 8.105653e-010,
  -3.592556e-013, 1.120659e-013, 7.173662e-011, 8.599806e-011,
  1.67623e-013, -7.693685e-016, -1.960875e-011, -7.806967e-011,
  5.028944e-014, 3.027491e-014, 1.046708e-010, 2.847257e-010,
  4.047984e-014, 7.635713e-014, 6.750647e-011, 5.6373e-011,
  9.157126e-014, 7.247545e-014, -5.823508e-011, -8.94328e-011,
  1.390933e-014, -3.567253e-014, -5.631789e-011, -1.313592e-010,
  -2.170292e-014, -2.889887e-014, 2.783449e-011, 3.1194e-011,
  -7.494832e-015, -3.451103e-014, 1.052868e-011, 2.636848e-011,
  -1.965583e-017, -8.342013e-015, 3.296329e-013, 2.682148e-012,
  -7.344484e-015, -6.155684e-014, -4.582281e-011, -9.413039e-011,
  9.389171e-015, -8.45247e-014, -5.083433e-012, 1.019504e-011,
  -2.862144e-013, 1.839373e-014, 6.213291e-011, 1.435064e-010,
  -1.456182e-014, 3.016655e-014, -1.608905e-010, -4.449902e-010,
  -1.413919e-013, -4.084271e-014, 5.683044e-011, 9.985431e-011,
  3.801156e-014, 8.888168e-014, -1.984745e-011, -1.107868e-010,
  6.943692e-014, -6.402841e-015, 4.045334e-011, 9.242392e-011,
  -3.42152e-014, -2.287349e-014, 6.663047e-011, 1.311617e-010,
  -1.689802e-013, 3.018295e-014, 1.877245e-010, 4.71747e-010,
  -1.852288e-013, 3.235093e-014, -8.637556e-011, -2.313891e-010,
  -9.843549e-014, 9.486626e-014, 7.70556e-011, 1.339441e-010,
  -3.527752e-014, 1.793312e-014, -1.260397e-010, -2.784702e-010,
  2.080624e-013, -9.115766e-014, -1.919723e-011, 4.580494e-011,
  -9.258579e-014, -1.329755e-014, 1.467004e-010, 3.272263e-010,
  3.223607e-013, -1.339854e-013, -3.42875e-010, -7.637204e-010,
  2.901871e-013, -1.622426e-013, 2.120834e-010, 5.534221e-010,
  1.057291e-012, -7.826678e-014, -4.603636e-010, -1.009472e-009,
  3.841396e-013, -3.279095e-013, 3.742011e-010, 1.152559e-009,
  -7.709553e-013, 4.291108e-014, -2.079138e-010, -5.293747e-010,
  4.658121e-013, -6.221132e-014, -5.427218e-010, -1.510281e-009,
  -2.066673e-014, 2.76431e-015, -1.010055e-010, -2.250616e-010,
  9.588808e-014, 6.577226e-014, 2.273904e-011, 3.734904e-011,
  1.758913e-013, -4.756508e-014, -1.768583e-011, 7.29451e-012,
  5.316376e-014, -4.131278e-014, 1.511264e-010, 4.580006e-010,
  3.81697e-013, 6.626259e-014, 5.537008e-010, 1.29478e-009,
  -8.021798e-013, 2.276716e-013, 1.747004e-010, 5.350733e-010,
  2.053955e-013, -1.022126e-013, 2.560653e-010, 5.775694e-010,
  -3.881474e-013, 2.933377e-014, 1.421327e-010, 4.013652e-010,
  -6.535282e-013, 9.722502e-014, 5.461851e-011, 2.521461e-010,
  -1.645997e-013, -1.080595e-013, -3.369504e-010, -9.263594e-010,
  -7.948795e-013, 1.624385e-013, 3.13885e-010, 7.672588e-010,
  -3.205715e-013, -1.118001e-014, -5.357806e-010, -1.305007e-009,
  -3.737079e-013, 1.754906e-014, -8.925177e-011, -1.437082e-010,
  1.592258e-013, -3.288211e-014, -2.022981e-010, -5.500759e-010,
  -4.950916e-013, 4.874728e-014, -1.38838e-011, 5.877309e-012,
  3.081356e-014, -2.764428e-014, -3.183309e-010, -8.516344e-010,
  4.874924e-013, -1.522703e-013, 1.170989e-010, 3.517102e-010,
  -2.881408e-013, 5.358615e-014, 4.030289e-010, 9.976914e-010,
  5.665406e-013, -1.489884e-013, 8.336477e-011, 2.355424e-010,
  -1.397352e-013, 1.42379e-014, 4.934971e-010, 1.231646e-009,
  -1.705243e-013, 4.133387e-014, 1.650965e-010, 4.348095e-010,
  -2.447336e-013, -1.089044e-014, -8.675603e-011, -2.456083e-010,
  -9.877415e-014, -7.431197e-014, 8.135266e-011, 2.183076e-010,
  -1.050358e-013, 4.064165e-015, 7.280729e-012, -1.259522e-011,
  -9.782665e-014, -1.234387e-014, 2.922913e-011, 7.363588e-011,
  1.888282e-014, 5.08231e-015, -5.903572e-011, -1.464635e-010,
  -2.872353e-013, -6.833604e-015, 3.539661e-010, 7.883426e-010,
  -1.665056e-013, 1.741338e-013, -1.389615e-010, -4.418301e-010,
  1.431109e-014, 1.540757e-014, -8.983745e-012, -4.095029e-011,
  -3.31204e-015, -2.986547e-014, -3.094792e-011, -4.248131e-011,
  -8.158357e-014, 2.387512e-014, 1.175736e-011, 3.669411e-011,
  7.757727e-015, -8.839083e-015, -9.100259e-011, -2.357962e-010,
  -1.062871e-012, 1.586071e-013, 6.261501e-010, 1.529722e-009,
  -6.771223e-013, 1.269877e-013, -5.35968e-010, -1.525654e-009,
  -1.071662e-013, -1.022993e-013, 3.407087e-010, 7.611797e-010,
  -2.693499e-013, 1.754659e-013, 1.328757e-010, 2.095504e-010,
  3.373075e-013, -5.919143e-014, 2.023801e-010, 2.172092e-010,
  6.501759e-014, 1.877695e-013, 2.835217e-010, 6.12537e-010,
  1.258924e-013, -1.162239e-013, -6.62818e-011, -1.84703e-010,
  2.047405e-014, 3.809218e-014, 1.588997e-010, 4.34363e-010,
  2.739003e-013, 3.454881e-013, 4.814769e-011, 1.523424e-010,
  -4.690994e-013, -2.179415e-013, -2.564357e-010, -4.705932e-010,
  -2.379047e-013, 1.039709e-013, 7.865346e-010, 1.987052e-009,
  -1.208172e-012, 2.272918e-013, 1.008904e-012, 3.666844e-011,
  8.732248e-014, -1.895771e-013, 1.334572e-010, 1.750704e-010,
  7.843009e-014, 1.730289e-013, 2.743864e-010, 5.57515e-010,
  4.676427e-013, 8.124497e-014, -8.585614e-011, 3.874778e-011,
  -2.372918e-013, 8.590089e-014, 2.89959e-010, 7.174599e-010,
  2.182818e-013, -9.436008e-014, 1.641019e-010, 2.974291e-010,
  -1.33482e-013, 2.02711e-013, 3.395071e-010, 7.9753e-010,
  -3.284387e-013, -1.763985e-013, 1.398132e-010, 3.17521e-010,
  -1.462416e-014, 1.26434e-013, 1.441746e-010, 6.397705e-011 ;

 emf_noise =
  3.537901e-015, 1.33519e-015, 2.072532e-011, 3.312415e-011,
  0, 0, 0, 0,
  6.740886e-015, 1.771798e-015, 2.66421e-011, 3.633482e-011,
  0, 0, 0, 0,
  1.821133e-014, 3.03556e-015, 3.687491e-011, 4.51221e-011,
  0, 0, 0, 0,
  6.845821e-014, 1.123475e-014, 5.63569e-011, 5.248878e-011,
  0, 0, 0, 0,
  1.313689e-014, 2.953949e-015, 3.017521e-011, 4.000054e-011,
  0, 0, 0, 0,
  7.440254e-015, 1.983686e-015, 3.279019e-011, 3.38444e-011,
  0, 0, 0, 0,
  5.450367e-014, 8.721039e-015, 4.71607e-011, 6.986218e-011,
  0, 0, 0, 0,
  5.638838e-015, 1.451898e-015, 2.326883e-011, 3.705393e-011,
  0, 0, 0, 0,
  5.775967e-015, 1.583676e-015, 2.96551e-011, 4.085247e-011,
  0, 0, 0, 0,
  1.997062e-014, 2.697061e-014, 1.866593e-011, 2.335805e-011,
  0, 0, 0, 0,
  5.173085e-014, 8.88147e-015, 2.316796e-011, 4.339543e-011,
  0, 0, 0, 0,
  1.087932e-014, 2.369893e-015, 2.438149e-011, 4.304743e-011,
  0, 0, 0, 0,
  8.065153e-014, 1.262482e-014, 3.166944e-011, 4.764645e-011,
  0, 0, 0, 0,
  1.086318e-014, 3.011139e-015, 3.981002e-011, 6.802179e-011,
  0, 0, 0, 0,
  6.325311e-015, 2.016338e-015, 2.495013e-011, 4.292542e-011,
  0, 0, 0, 0,
  1.324001e-014, 3.300167e-015, 2.987195e-011, 6.291916e-011,
  0, 0, 0, 0,
  2.949497e-014, 5.448606e-015, 6.863594e-011, 1.164782e-010,
  0, 0, 0, 0,
  1.042943e-014, 2.013209e-015, 1.59719e-011, 3.46982e-011,
  0, 0, 0, 0,
  1.111316e-014, 2.872675e-015, 1.769749e-011, 2.739743e-011,
  0, 0, 0, 0,
  7.477791e-015, 2.752894e-015, 1.890316e-011, 2.49088e-011,
  0, 0, 0, 0,
  9.238359e-015, 2.635359e-015, 3.883094e-011, 6.108188e-011,
  0, 0, 0, 0,
  7.573062e-015, 1.823797e-015, 2.549676e-011, 3.99426e-011,
  0, 0, 0, 0,
  1.364774e-014, 3.089397e-015, 4.304548e-011, 7.312525e-011,
  0, 0, 0, 0,
  6.457831e-014, 1.054206e-014, 4.882426e-011, 7.780784e-011,
  0, 0, 0, 0,
  1.648367e-014, 5.341392e-015, 3.623895e-011, 5.985872e-011,
  0, 0, 0, 0,
  1.840323e-014, 3.972115e-015, 3.777651e-011, 5.383833e-011,
  0, 0, 0, 0,
  2.414928e-014, 4.021266e-015, 3.543649e-011, 6.353566e-011,
  0, 0, 0, 0,
  5.512379e-014, 8.802729e-015, 5.897345e-011, 8.416641e-011,
  0, 0, 0, 0,
  2.664784e-014, 5.65579e-015, 4.246889e-011, 6.560023e-011,
  0, 0, 0, 0,
  3.78368e-014, 6.234623e-015, 5.303783e-011, 7.307946e-011,
  0, 0, 0, 0,
  7.099205e-015, 1.581492e-015, 1.32168e-011, 2.349311e-011,
  0, 0, 0, 0,
  7.818477e-015, 1.737695e-015, 2.42065e-011, 4.700538e-011,
  0, 0, 0, 0,
  1.774807e-014, 3.381371e-015, 5.532207e-011, 9.980437e-011,
  0, 0, 0, 0,
  1.031647e-014, 2.086201e-015, 1.988072e-011, 3.465263e-011,
  0, 0, 0, 0,
  3.031216e-014, 5.008331e-015, 3.585907e-011, 5.912723e-011,
  0, 0, 0, 0,
  3.952042e-014, 6.6017e-015, 4.238547e-011, 6.005085e-011,
  0, 0, 0, 0,
  2.485757e-014, 4.664552e-015, 4.087068e-011, 6.173281e-011,
  0, 0, 0, 0,
  2.289272e-014, 4.151697e-015, 3.443495e-011, 4.735717e-011,
  0, 0, 0, 0,
  7.479259e-015, 1.569759e-015, 2.195602e-011, 3.475329e-011,
  0, 0, 0, 0,
  1.487289e-014, 2.582106e-015, 2.462533e-011, 3.438074e-011,
  0, 0, 0, 0,
  4.586076e-014, 7.302501e-015, 3.321932e-011, 5.209448e-011,
  0, 0, 0, 0,
  8.20674e-015, 2.255466e-015, 3.604752e-011, 5.923963e-011,
  0, 0, 0, 0,
  5.835501e-015, 1.754215e-015, 2.99443e-011, 4.288258e-011,
  0, 0, 0, 0,
  4.607096e-015, 2.322718e-015, 5.287146e-011, 7.814138e-011,
  0, 0, 0, 0,
  5.908979e-014, 9.122634e-015, 1.382029e-011, 2.234846e-011,
  0, 0, 0, 0,
  2.194362e-014, 3.89393e-015, 3.206801e-011, 2.692534e-011,
  0, 0, 0, 0,
  1.852405e-014, 3.958576e-015, 2.257247e-011, 2.271971e-011,
  0, 0, 0, 0,
  1.8848e-014, 3.224127e-015, 1.880399e-011, 2.148921e-011,
  0, 0, 0, 0,
  3.878421e-014, 1.732673e-014, 1.909751e-011, 2.643315e-011,
  0, 0, 0, 0,
  2.618312e-014, 4.499342e-015, 1.905233e-011, 1.467676e-011,
  0, 0, 0, 0,
  2.11179e-014, 4.572233e-015, 1.324251e-011, 3.159476e-011,
  0, 0, 0, 0,
  3.201652e-014, 5.440035e-015, 8.309645e-012, 1.421132e-011,
  0, 0, 0, 0,
  4.349657e-014, 7.293645e-015, 2.068602e-011, 3.104127e-011,
  0, 0, 0, 0,
  4.854171e-014, 8.261266e-015, 2.302554e-011, 3.346142e-011,
  0, 0, 0, 0,
  1.037065e-014, 2.031817e-015, 2.644377e-011, 3.792803e-011,
  0, 0, 0, 0,
  1.511987e-014, 3.157487e-015, 4.184171e-011, 5.469379e-011,
  0, 0, 0, 0,
  1.753877e-014, 2.84792e-015, 2.153078e-011, 3.545069e-011,
  0, 0, 0, 0,
  4.361515e-014, 6.935422e-015, 4.697581e-011, 7.72277e-011,
  0, 0, 0, 0,
  2.062761e-014, 4.061857e-015, 2.94761e-011, 3.490932e-011,
  0, 0, 0, 0,
  1.348339e-014, 2.302718e-015, 7.979321e-012, 1.014128e-011,
  0, 0, 0, 0,
  2.383098e-014, 4.266718e-015, 9.701641e-012, 1.408595e-011,
  0, 0, 0, 0,
  1.198113e-014, 2.273751e-015, 1.295993e-011, 2.173608e-011,
  0, 0, 0, 0,
  7.048031e-015, 2.017117e-015, 1.615158e-011, 2.764321e-011,
  0, 0, 0, 0,
  1.671695e-014, 2.690568e-015, 9.903262e-012, 8.574486e-012,
  0, 0, 0, 0,
  7.954653e-015, 1.732623e-015, 9.704343e-012, 1.639129e-011,
  0, 0, 0, 0,
  3.158559e-014, 5.392863e-015, 2.310277e-011, 2.119428e-011,
  0, 0, 0, 0,
  1.139445e-014, 3.205976e-015, 2.560062e-011, 3.76266e-011,
  0, 0, 0, 0,
  2.068911e-014, 4.08551e-015, 3.499997e-011, 3.854671e-011,
  0, 0, 0, 0,
  5.616068e-014, 9.339682e-015, 6.349494e-011, 9.235609e-011,
  0, 0, 0, 0,
  4.512633e-014, 7.413639e-015, 3.328037e-011, 4.645178e-011,
  0, 0, 0, 0,
  1.33498e-014, 2.670406e-015, 3.200636e-011, 5.297922e-011,
  0, 0, 0, 0,
  9.438564e-015, 2.064065e-015, 2.986997e-011, 3.468175e-011,
  0, 0, 0, 0,
  7.558858e-015, 2.28669e-015, 2.590508e-011, 3.914326e-011,
  0, 0, 0, 0,
  2.757342e-014, 4.606432e-015, 1.193437e-011, 1.675005e-011,
  0, 0, 0, 0,
  4.162524e-014, 6.441719e-015, 2.347087e-011, 3.730108e-011,
  0, 0, 0, 0,
  1.941106e-014, 3.526807e-015, 3.017313e-011, 4.038323e-011,
  0, 0, 0, 0,
  1.353105e-014, 2.650021e-015, 1.845384e-011, 2.487047e-011,
  0, 0, 0, 0,
  1.011348e-014, 2.700028e-015, 2.162467e-011, 3.072561e-011,
  0, 0, 0, 0,
  3.426979e-014, 5.885601e-015, 6.260731e-011, 6.656441e-011,
  0, 0, 0, 0,
  2.580714e-014, 4.781117e-015, 7.000087e-011, 7.925158e-011,
  0, 0, 0, 0,
  1.23486e-014, 3.176078e-015, 7.159753e-011, 9.922579e-011,
  0, 0, 0, 0,
  2.990263e-014, 6.26069e-015, 1.162581e-010, 1.449229e-010,
  0, 0, 0, 0,
  1.332143e-014, 3.276365e-015, 5.370429e-011, 6.49317e-011,
  0, 0, 0, 0,
  1.333584e-014, 3.312483e-015, 7.566143e-011, 7.863293e-011,
  0, 0, 0, 0,
  9.285511e-015, 3.020383e-015, 7.701835e-011, 8.890702e-011,
  0, 0, 0, 0,
  8.832085e-015, 4.770466e-015, 7.254804e-011, 1.00618e-010,
  0, 0, 0, 0,
  5.483318e-014, 8.717959e-015, 2.041389e-011, 2.223875e-011,
  0, 0, 0, 0,
  9.317346e-015, 3.523614e-015, 2.507521e-011, 3.281947e-011,
  0, 0, 0, 0,
  8.357801e-015, 2.267551e-015, 2.716394e-011, 2.303237e-011,
  0, 0, 0, 0,
  3.069296e-014, 6.278266e-015, 1.219404e-010, 1.230799e-010,
  0, 0, 0, 0,
  3.680547e-014, 6.130545e-015, 6.404088e-011, 5.702036e-011,
  0, 0, 0, 0,
  2.101518e-014, 3.561833e-015, 3.018272e-011, 2.979614e-011,
  0, 0, 0, 0,
  1.283413e-014, 3.929737e-015, 5.966231e-011, 6.154637e-011,
  0, 0, 0, 0,
  1.269189e-014, 2.958802e-015, 5.957157e-011, 7.470546e-011,
  0, 0, 0, 0,
  2.236106e-014, 4.205348e-015, 5.030633e-011, 5.602501e-011,
  0, 0, 0, 0,
  1.848608e-014, 4.358755e-015, 4.574407e-011, 4.81092e-011,
  0, 0, 0, 0,
  6.211931e-015, 4.40761e-015, 4.695475e-011, 6.426519e-011,
  0, 0, 0, 0,
  1.422606e-014, 4.605031e-015, 2.773004e-011, 4.561792e-011,
  0, 0, 0, 0,
  1.955429e-014, 5.467783e-015, 4.591076e-011, 6.213051e-011,
  0, 0, 0, 0,
  1.632917e-014, 3.462656e-015, 1.69218e-011, 1.255671e-011,
  0, 0, 0, 0,
  8.467133e-015, 3.24034e-015, 1.135741e-011, 1.414937e-011,
  0, 0, 0, 0,
  5.348866e-015, 3.338338e-015, 1.411943e-011, 1.41928e-011,
  0, 0, 0, 0,
  1.029943e-014, 4.544272e-015, 2.145786e-011, 2.622654e-011,
  0, 0, 0, 0,
  1.662842e-014, 4.761808e-015, 3.808973e-011, 4.333691e-011,
  0, 0, 0, 0,
  1.031059e-014, 3.569162e-015, 5.293967e-011, 6.524636e-011,
  0, 0, 0, 0,
  2.393184e-014, 6.461127e-015, 7.06122e-011, 8.771315e-011,
  0, 0, 0, 0,
  1.12394e-014, 4.668059e-015, 2.291528e-011, 2.398627e-011,
  0, 0, 0, 0,
  1.838006e-014, 5.44589e-015, 8.154233e-011, 8.230003e-011,
  0, 0, 0, 0,
  1.790347e-014, 1.428886e-014, 1.840991e-010, 2.076056e-010,
  0, 0, 0, 0,
  1.148686e-014, 6.957484e-015, 4.186685e-011, 3.641181e-011,
  0, 0, 0, 0,
  1.807313e-014, 7.887829e-015, 5.506539e-011, 6.979019e-011,
  0, 0, 0, 0,
  1.828909e-014, 7.338897e-015, 2.194017e-011, 1.707038e-011,
  0, 0, 0, 0,
  2.318651e-014, 1.107418e-014, 1.46453e-011, 1.476874e-011,
  0, 0, 0, 0,
  3.364413e-014, 8.871373e-015, 2.182264e-011, 3.615546e-011,
  0, 0, 0, 0,
  3.983304e-014, 1.100544e-014, 2.399542e-011, 2.778689e-011,
  0, 0, 0, 0,
  6.085283e-014, 1.245258e-014, 3.031492e-011, 2.468841e-011,
  0, 0, 0, 0,
  5.149955e-014, 1.423264e-014, 3.164683e-011, 3.767119e-011,
  0, 0, 0, 0,
  6.966636e-014, 1.924613e-014, 4.513806e-011, 5.427764e-011,
  0, 0, 0, 0,
  7.514435e-014, 4.929146e-014, 2.684019e-011, 2.643607e-011,
  0, 0, 0, 0,
  1.072012e-012, 1.769746e-013, 3.432817e-011, 6.529163e-011,
  0, 0, 0, 0,
  1.567836e-013, 5.341052e-014, 2.403377e-011, 3.071235e-011,
  0, 0, 0, 0,
  2.112023e-013, 5.605953e-014, 5.522386e-011, 5.267103e-011,
  0, 0, 0, 0,
  3.336805e-013, 8.621993e-014, 4.967006e-011, 5.573529e-011,
  0, 0, 0, 0,
  5.458349e-013, 1.397872e-013, 4.219914e-011, 9.266202e-011,
  0, 0, 0, 0,
  9.02447e-013, 2.128593e-013, 1.188752e-010, 3.067221e-010,
  0, 0, 0, 0,
  1.530379e-012, 4.362529e-013, 1.629496e-010, 3.295175e-010,
  0, 0, 0, 0,
  2.333575e-012, 7.17101e-013, 3.362859e-010, 5.306914e-010,
  0, 0, 0, 0,
  3.266288e-012, 2.041683e-012, 5.716025e-010, 1.348329e-009,
  0, 0, 0, 0,
  1.283403e-011, 3.479936e-012, 1.180067e-009, 6.21127e-009,
  0, 0, 0, 0,
  1.060218e-011, 3.486133e-012, 5.761807e-010, 1.614482e-009,
  0, 0, 0, 0,
  2.674441e-012, 1.677483e-012, 4.395872e-010, 7.730491e-010,
  0, 0, 0, 0,
  1.161131e-011, 2.76248e-012, 6.775479e-010, 1.947753e-009,
  0, 0, 0, 0,
  1.171875e-011, 3.472565e-012, 5.852507e-010, 1.966063e-009,
  0, 0, 0, 0,
  2.782001e-012, 2.06687e-012, 3.077692e-010, 1.107511e-009,
  0, 0, 0, 0,
  2.403279e-012, 5.116099e-013, 1.433427e-010, 4.664265e-010,
  0, 0, 0, 0,
  1.474901e-012, 4.060523e-013, 6.97872e-011, 2.292381e-010,
  0, 0, 0, 0,
  7.741772e-013, 2.564872e-013, 4.025406e-011, 1.260138e-010,
  0, 0, 0, 0,
  4.776066e-013, 1.756783e-013, 5.082016e-011, 8.639552e-011,
  0, 0, 0, 0,
  3.295322e-013, 9.757078e-014, 6.065392e-011, 7.465065e-011,
  0, 0, 0, 0,
  2.308237e-013, 5.696241e-014, 3.036675e-011, 4.061785e-011,
  0, 0, 0, 0,
  1.555985e-013, 6.536839e-014, 3.039449e-011, 3.179198e-011,
  0, 0, 0, 0,
  1.082677e-013, 4.872692e-014, 2.802097e-011, 4.649917e-011,
  0, 0, 0, 0,
  8.735809e-014, 2.196223e-014, 4.291498e-011, 3.296109e-011,
  0, 0, 0, 0,
  6.136127e-014, 1.833316e-014, 3.886995e-011, 3.921333e-011,
  0, 0, 0, 0,
  5.829152e-014, 1.74731e-014, 4.441053e-011, 4.85464e-011,
  0, 0, 0, 0,
  5.16787e-014, 1.291092e-014, 2.666546e-011, 2.688001e-011,
  0, 0, 0, 0,
  3.555084e-014, 1.356109e-014, 1.058965e-011, 1.419639e-011,
  0, 0, 0, 0,
  2.637153e-014, 8.200212e-015, 1.551009e-011, 2.541403e-011,
  0, 0, 0, 0,
  2.469781e-014, 1.299708e-014, 1.10185e-011, 1.76056e-011,
  0, 0, 0, 0,
  2.19681e-014, 4.929917e-015, 2.146935e-011, 2.758731e-011,
  0, 0, 0, 0,
  2.790168e-014, 1.160859e-014, 2.982115e-011, 6.100505e-011,
  0, 0, 0, 0,
  1.341205e-014, 7.649403e-015, 3.612707e-011, 5.563135e-011,
  0, 0, 0, 0,
  1.265584e-014, 5.243272e-015, 4.276232e-011, 1.037374e-010,
  0, 0, 0, 0,
  5.409239e-014, 2.552483e-014, 5.253687e-011, 4.415582e-011,
  0, 0, 0, 0,
  1.263377e-014, 1.033745e-014, 2.665772e-011, 5.714755e-011,
  0, 0, 0, 0,
  6.475813e-015, 8.445363e-015, 4.313126e-011, 8.66431e-011,
  0, 0, 0, 0,
  6.699554e-015, 3.269339e-015, 1.817227e-011, 2.595486e-011,
  0, 0, 0, 0,
  5.62923e-015, 2.881638e-015, 2.847052e-011, 1.674672e-011,
  0, 0, 0, 0,
  7.443283e-015, 3.650343e-015, 2.555818e-011, 3.608589e-011,
  0, 0, 0, 0,
  5.790962e-015, 4.290747e-015, 4.780373e-011, 5.17489e-011,
  0, 0, 0, 0,
  4.746912e-015, 3.339315e-015, 2.701319e-011, 2.262626e-011,
  0, 0, 0, 0,
  4.55047e-015, 6.361504e-015, 6.665308e-011, 3.332117e-011,
  0, 0, 0, 0,
  4.982711e-015, 5.646831e-015, 3.128564e-011, 3.897433e-011,
  0, 0, 0, 0,
  2.895917e-015, 3.070632e-015, 2.010582e-011, 1.935309e-011,
  0, 0, 0, 0,
  4.012249e-015, 4.574487e-015, 2.768284e-011, 2.871237e-011,
  0, 0, 0, 0,
  1.974109e-015, 1.942204e-015, 1.865778e-011, 1.696064e-011,
  0, 0, 0, 0,
  2.650817e-015, 1.77301e-015, 1.440422e-011, 1.238627e-011,
  0, 0, 0, 0,
  2.578979e-015, 4.674873e-015, 2.644779e-011, 2.040218e-011,
  0, 0, 0, 0,
  4.680706e-015, 3.028714e-015, 2.887682e-011, 5.851686e-011,
  0, 0, 0, 0,
  4.324279e-015, 6.249344e-015, 4.447006e-011, 1.907569e-011,
  0, 0, 0, 0,
  9.963857e-015, 3.130448e-015, 1.992995e-011, 2.957111e-011,
  0, 0, 0, 0,
  3.548573e-015, 6.325213e-015, 5.017812e-011, 6.215137e-011,
  0, 0, 0, 0,
  3.407607e-015, 5.122024e-015, 3.437825e-011, 4.956395e-011,
  0, 0, 0, 0,
  2.285066e-015, 2.889705e-015, 1.988734e-011, 2.217949e-011,
  0, 0, 0, 0,
  4.78579e-014, 8.009577e-015, 2.718929e-011, 1.932355e-011,
  0, 0, 0, 0,
  8.151229e-015, 4.424901e-015, 4.271225e-011, 3.363093e-011,
  0, 0, 0, 0,
  2.208816e-015, 2.632059e-015, 2.240848e-011, 1.723425e-011,
  0, 0, 0, 0,
  1.803013e-015, 7.251818e-015, 3.097773e-011, 2.4342e-011,
  0, 0, 0, 0,
  3.383523e-014, 7.227624e-015, 5.905453e-011, 4.447415e-011,
  0, 0, 0, 0,
  2.134218e-014, 3.869154e-015, 1.623457e-011, 1.57285e-011,
  0, 0, 0, 0,
  5.677994e-015, 4.32846e-015, 4.847575e-011, 2.917668e-011,
  0, 0, 0, 0,
  4.040508e-015, 4.621405e-015, 4.637528e-011, 5.779322e-011,
  0, 0, 0, 0,
  4.310189e-015, 5.555115e-015, 7.538618e-011, 5.675319e-011,
  0, 0, 0, 0,
  3.964828e-015, 3.425709e-015, 3.557193e-011, 6.145292e-011,
  0, 0, 0, 0,
  1.822779e-015, 7.787551e-015, 6.403197e-011, 4.495442e-011,
  0, 0, 0, 0,
  2.889068e-015, 4.94476e-015, 2.534812e-011, 5.827991e-011,
  0, 0, 0, 0,
  3.052289e-015, 7.013457e-015, 3.693209e-011, 3.52698e-011,
  0, 0, 0, 0,
  7.299915e-015, 4.131204e-015, 1.777094e-011, 1.715913e-011,
  0, 0, 0, 0,
  3.063518e-015, 7.204243e-015, 5.61528e-011, 3.778184e-011,
  0, 0, 0, 0,
  5.452002e-015, 7.895812e-015, 3.218332e-011, 6.780851e-011,
  0, 0, 0, 0,
  3.222719e-015, 4.959839e-015, 2.866687e-011, 3.511217e-011,
  0, 0, 0, 0,
  4.973352e-014, 7.792104e-015, 1.033132e-011, 9.024527e-012,
  0, 0, 0, 0,
  2.541176e-015, 2.499191e-015, 1.963274e-011, 2.766067e-011,
  0, 0, 0, 0,
  3.95943e-015, 2.658124e-015, 3.490671e-011, 2.226643e-011,
  0, 0, 0, 0,
  2.439303e-015, 2.802426e-015, 2.880688e-011, 2.126932e-011,
  0, 0, 0, 0,
  4.079291e-014, 6.55304e-015, 1.832344e-011, 1.072122e-011,
  0, 0, 0, 0,
  1.357891e-014, 3.334663e-015, 1.563784e-011, 2.997645e-011,
  0, 0, 0, 0,
  2.12435e-015, 2.488411e-015, 2.063764e-011, 1.910952e-011,
  0, 0, 0, 0,
  1.103335e-015, 3.283609e-015, 2.345336e-011, 1.654774e-011,
  0, 0, 0, 0,
  1.614876e-015, 3.386834e-015, 3.504465e-011, 3.111789e-011,
  0, 0, 0, 0,
  7.959645e-016, 3.896693e-015, 4.054532e-011, 2.936355e-011,
  0, 0, 0, 0,
  2.133364e-015, 2.512361e-015, 1.761103e-011, 2.480507e-011,
  0, 0, 0, 0,
  1.479226e-015, 3.58941e-015, 4.163964e-011, 2.687894e-011,
  0, 0, 0, 0,
  1.997959e-015, 1.76802e-015, 2.014422e-011, 3.568436e-011,
  0, 0, 0, 0,
  5.662323e-015, 3.732923e-015, 2.796743e-011, 4.343151e-011,
  0, 0, 0, 0,
  2.03926e-015, 2.571685e-015, 3.459829e-011, 2.631342e-011,
  0, 0, 0, 0,
  2.809849e-015, 6.343716e-015, 6.358596e-011, 8.265508e-011,
  0, 0, 0, 0,
  3.360164e-015, 4.95366e-015, 5.26043e-011, 9.945463e-011,
  0, 0, 0, 0,
  5.108435e-014, 8.898535e-015, 3.384176e-011, 4.706627e-011,
  0, 0, 0, 0,
  4.370529e-015, 5.567191e-015, 3.475568e-011, 4.300839e-011,
  0, 0, 0, 0,
  5.523954e-015, 1.612975e-014, 4.128513e-011, 6.910066e-011,
  0, 0, 0, 0,
  1.899709e-015, 1.629759e-015, 3.214375e-011, 4.073425e-011,
  0, 0, 0, 0,
  4.557866e-014, 7.616123e-015, 3.943644e-011, 5.130494e-011,
  0, 0, 0, 0,
  9.210141e-015, 3.115424e-015, 2.980434e-011, 2.818521e-011,
  0, 0, 0, 0,
  2.771352e-015, 2.39268e-015, 3.115213e-011, 3.960623e-011,
  0, 0, 0, 0,
  3.081301e-015, 4.166727e-015, 3.273392e-011, 4.03898e-011,
  0, 0, 0, 0,
  5.204912e-015, 4.31929e-015, 4.111795e-011, 6.931182e-011,
  0, 0, 0, 0,
  3.786178e-015, 2.796431e-015, 6.185065e-011, 7.464891e-011,
  0, 0, 0, 0,
  5.590776e-015, 4.695553e-015, 7.292151e-011, 8.519187e-011,
  0, 0, 0, 0,
  2.759408e-015, 5.783257e-015, 3.048454e-011, 4.603786e-011,
  0, 0, 0, 0,
  1.686072e-014, 5.086941e-015, 3.005075e-011, 4.386116e-011,
  0, 0, 0, 0,
  3.865893e-014, 6.260697e-015, 4.281317e-011, 4.596456e-011,
  0, 0, 0, 0,
  2.059914e-015, 2.950785e-015, 2.935257e-011, 5.449456e-011,
  0, 0, 0, 0,
  1.686735e-015, 2.12518e-015, 1.65829e-011, 2.064531e-011,
  0, 0, 0, 0,
  3.08927e-015, 1.984631e-015, 2.309325e-011, 4.267942e-011,
  0, 0, 0, 0,
  5.448924e-014, 9.073079e-015, 5.512519e-011, 5.031305e-011,
  0, 0, 0, 0,
  2.780131e-015, 2.203746e-015, 4.141325e-011, 6.66621e-011,
  0, 0, 0, 0,
  4.844617e-015, 2.811324e-015, 3.749448e-011, 5.566369e-011,
  0, 0, 0, 0,
  4.588234e-015, 3.168022e-015, 2.100336e-011, 5.789682e-011,
  0, 0, 0, 0,
  3.716675e-015, 3.289655e-015, 1.667609e-011, 2.024976e-011,
  0, 0, 0, 0,
  1.6909e-015, 3.288484e-015, 1.544919e-011, 2.478804e-011,
  0, 0, 0, 0,
  1.126307e-015, 2.180982e-015, 8.495929e-012, 1.87749e-011,
  0, 0, 0, 0,
  9.061003e-015, 3.565213e-015, 1.326225e-011, 3.795756e-011,
  0, 0, 0, 0,
  3.742955e-014, 6.029349e-015, 3.233526e-011, 5.480803e-011,
  0, 0, 0, 0,
  1.797621e-014, 3.370457e-015, 2.04695e-011, 1.387031e-011,
  0, 0, 0, 0,
  5.070262e-014, 8.125962e-015, 4.0612e-011, 3.266187e-011,
  0, 0, 0, 0,
  1.12801e-014, 3.997739e-015, 3.596086e-011, 6.818979e-011,
  0, 0, 0, 0,
  1.903457e-014, 3.608314e-015, 2.135157e-011, 4.491056e-011,
  0, 0, 0, 0,
  3.808701e-014, 6.37122e-015, 1.977178e-011, 4.00435e-011,
  0, 0, 0, 0,
  2.912547e-015, 2.452044e-015, 2.164797e-011, 3.762483e-011,
  0, 0, 0, 0,
  2.775254e-015, 1.996057e-015, 2.208658e-011, 5.80726e-011,
  0, 0, 0, 0,
  1.495475e-015, 3.081886e-015, 1.236353e-011, 2.085465e-011,
  0, 0, 0, 0,
  3.151406e-015, 2.233078e-015, 4.546935e-011, 5.357422e-011,
  0, 0, 0, 0,
  2.357263e-015, 2.823979e-015, 2.264669e-011, 2.82258e-011,
  0, 0, 0, 0,
  2.302185e-015, 1.366492e-015, 2.01231e-011, 3.037127e-011,
  0, 0, 0, 0,
  2.554683e-015, 2.628308e-015, 1.426096e-011, 3.120885e-011,
  0, 0, 0, 0,
  5.135583e-014, 8.221967e-015, 2.381499e-011, 1.886947e-011,
  0, 0, 0, 0,
  2.078023e-015, 2.461669e-015, 2.463149e-011, 3.198975e-011,
  0, 0, 0, 0,
  3.291141e-015, 3.602144e-015, 2.121477e-011, 5.100788e-011,
  0, 0, 0, 0,
  4.010465e-015, 2.891944e-015, 2.10499e-011, 3.277467e-011,
  0, 0, 0, 0,
  4.269179e-014, 7.055311e-015, 4.246272e-011, 9.943662e-011,
  0, 0, 0, 0,
  1.471913e-014, 6.806504e-015, 3.430174e-011, 5.185148e-011,
  0, 0, 0, 0,
  2.258953e-015, 3.497387e-015, 3.802558e-011, 5.642039e-011,
  0, 0, 0, 0,
  4.376275e-015, 5.567496e-015, 4.531238e-011, 4.041688e-011,
  0, 0, 0, 0,
  4.135599e-015, 4.078946e-015, 4.031938e-011, 4.950396e-011,
  0, 0, 0, 0,
  2.922907e-015, 4.106953e-015, 3.552008e-011, 4.533766e-011,
  0, 0, 0, 0,
  4.102415e-015, 4.408378e-015, 3.610267e-011, 6.298961e-011,
  0, 0, 0, 0,
  1.922828e-015, 3.045467e-015, 3.654322e-011, 5.068427e-011,
  0, 0, 0, 0,
  8.750166e-015, 2.701211e-015, 3.54701e-011, 8.070387e-011,
  0, 0, 0, 0,
  4.698547e-014, 7.360551e-015, 1.202637e-011, 1.361635e-011,
  0, 0, 0, 0,
  1.975247e-015, 1.444641e-015, 2.680347e-011, 3.106954e-011,
  0, 0, 0, 0,
  2.2477e-015, 1.283906e-015, 2.952187e-011, 2.409704e-011,
  0, 0, 0, 0,
  1.765672e-015, 1.776817e-015, 1.856375e-011, 2.091019e-011,
  0, 0, 0, 0,
  5.484051e-014, 8.639944e-015, 2.095519e-011, 3.180661e-011,
  0, 0, 0, 0,
  2.044902e-015, 2.317867e-015, 1.624485e-011, 1.590415e-011,
  0, 0, 0, 0,
  2.819307e-015, 2.391804e-015, 3.954049e-011, 2.747618e-011,
  0, 0, 0, 0,
  5.180222e-015, 4.95857e-015, 3.708659e-011, 6.038228e-011,
  0, 0, 0, 0,
  2.848019e-015, 2.382922e-015, 4.459135e-011, 8.258588e-011,
  0, 0, 0, 0,
  2.76802e-015, 2.483506e-015, 2.608975e-011, 3.144475e-011,
  0, 0, 0, 0,
  2.07964e-015, 2.854531e-015, 2.694993e-011, 3.999312e-011,
  0, 0, 0, 0,
  2.069744e-015, 4.569911e-015, 3.588954e-011, 7.282943e-011,
  0, 0, 0, 0,
  2.559716e-015, 2.852496e-015, 2.520959e-011, 4.034006e-011,
  0, 0, 0, 0,
  4.976994e-015, 2.531191e-015, 2.450165e-011, 2.640301e-011,
  0, 0, 0, 0,
  3.247715e-015, 4.177128e-015, 3.462048e-011, 4.437457e-011,
  0, 0, 0, 0,
  2.218751e-015, 5.164445e-015, 2.027977e-011, 3.7442e-011,
  0, 0, 0, 0,
  1.386487e-014, 4.351493e-015, 2.426153e-011, 3.671458e-011,
  0, 0, 0, 0,
  4.059402e-014, 8.025077e-015, 3.029283e-011, 4.864604e-011,
  0, 0, 0, 0,
  1.899411e-015, 3.697123e-015, 4.067663e-011, 4.661212e-011,
  0, 0, 0, 0,
  3.168934e-015, 2.523744e-015, 2.117904e-011, 3.116206e-011,
  0, 0, 0, 0,
  2.306129e-015, 3.652292e-015, 2.189119e-011, 2.598654e-011,
  0, 0, 0, 0,
  5.182235e-014, 8.284918e-015, 9.371098e-012, 1.213234e-011,
  0, 0, 0, 0,
  2.325019e-015, 1.859689e-015, 1.223585e-011, 2.32959e-011,
  0, 0, 0, 0,
  3.670099e-015, 3.357208e-015, 2.712192e-011, 5.678244e-011,
  0, 0, 0, 0,
  3.151403e-015, 3.222546e-015, 2.800697e-011, 4.968833e-011,
  0, 0, 0, 0,
  2.64319e-015, 3.363343e-015, 2.494959e-011, 4.204184e-011,
  0, 0, 0, 0,
  2.504474e-015, 4.403435e-015, 2.901106e-011, 3.804998e-011,
  0, 0, 0, 0,
  1.890052e-015, 2.922313e-015, 1.027328e-011, 1.992208e-011,
  0, 0, 0, 0,
  1.493606e-015, 1.954672e-015, 1.718568e-011, 2.507783e-011,
  0, 0, 0, 0,
  4.312879e-014, 7.206264e-015, 1.794175e-011, 3.48497e-011,
  0, 0, 0, 0,
  1.339857e-014, 4.111575e-015, 2.6663e-011, 3.256452e-011,
  0, 0, 0, 0,
  5.292795e-015, 3.030432e-015, 4.464188e-011, 6.374e-011,
  0, 0, 0, 0,
  4.1029e-015, 3.794358e-015, 3.889842e-011, 5.222496e-011,
  0, 0, 0, 0,
  2.250249e-014, 4.619099e-015, 3.580761e-011, 4.665853e-011,
  0, 0, 0, 0,
  3.954357e-014, 7.522129e-015, 3.591063e-011, 6.184012e-011,
  0, 0, 0, 0,
  3.937832e-015, 4.880201e-015, 3.855655e-011, 6.341434e-011,
  0, 0, 0, 0,
  3.934727e-015, 3.749602e-015, 5.897319e-011, 8.866134e-011,
  0, 0, 0, 0,
  1.743822e-015, 2.793446e-015, 3.590869e-011, 7.779521e-011,
  0, 0, 0, 0,
  1.827171e-015, 2.232119e-015, 1.759195e-011, 2.749147e-011,
  0, 0, 0, 0,
  2.704385e-015, 3.171028e-015, 1.687593e-011, 4.6578e-011,
  0, 0, 0, 0,
  2.257302e-015, 3.496681e-015, 2.202157e-011, 5.44646e-011,
  0, 0, 0, 0,
  3.054272e-015, 2.595746e-015, 2.946343e-011, 5.182883e-011,
  0, 0, 0, 0,
  5.070743e-014, 8.441535e-015, 2.440412e-011, 4.621618e-011,
  0, 0, 0, 0,
  1.843515e-015, 1.444902e-015, 2.225122e-011, 2.095397e-011,
  0, 0, 0, 0,
  3.20473e-015, 2.165699e-015, 2.468091e-011, 3.295737e-011,
  0, 0, 0, 0,
  1.526694e-015, 2.651319e-015, 2.124099e-011, 2.884337e-011,
  0, 0, 0, 0,
  4.632361e-014, 7.384281e-015, 2.477339e-011, 4.883868e-011,
  0, 0, 0, 0,
  9.313425e-015, 2.529759e-015, 1.783403e-011, 3.078171e-011,
  0, 0, 0, 0,
  2.955091e-015, 2.053709e-015, 3.005312e-011, 5.570174e-011,
  0, 0, 0, 0,
  1.496162e-015, 1.98617e-015, 1.814108e-011, 1.652519e-011,
  0, 0, 0, 0,
  2.216882e-015, 3.516637e-015, 2.047177e-011, 1.670547e-011,
  0, 0, 0, 0,
  2.730596e-015, 4.539046e-015, 2.129825e-011, 4.010228e-011,
  0, 0, 0, 0,
  5.486805e-015, 2.793737e-015, 3.275392e-011, 5.21086e-011,
  0, 0, 0, 0,
  3.201984e-015, 5.120221e-015, 4.804436e-011, 1.036154e-010,
  0, 0, 0, 0,
  2.72321e-015, 3.138374e-015, 4.227977e-011, 6.381992e-011,
  0, 0, 0, 0,
  6.189911e-015, 3.172268e-015, 3.096051e-011, 5.151492e-011,
  0, 0, 0, 0,
  3.763713e-015, 3.967332e-015, 8.07774e-011, 1.374355e-010,
  0, 0, 0, 0,
  3.651876e-015, 3.225878e-015, 3.77235e-011, 6.534695e-011,
  0, 0, 0, 0,
  5.285642e-015, 5.237147e-015, 7.420788e-011, 8.3373e-011,
  0, 0, 0, 0,
  1.466671e-015, 1.945352e-015, 3.508057e-012, 5.083236e-012,
  0, 0, 0, 0,
  6.165587e-015, 2.040542e-015, 1.773567e-011, 1.082752e-011,
  0, 0, 0, 0,
  2.54177e-014, 4.774604e-015, 6.815518e-012, 1.025472e-011,
  0, 0, 0, 0,
  3.338854e-014, 6.045758e-015, 2.572012e-011, 3.028688e-011,
  0, 0, 0, 0,
  4.03475e-015, 2.846154e-015, 7.506185e-012, 1.195465e-011,
  0, 0, 0, 0,
  1.218697e-015, 2.445102e-015, 9.396229e-012, 9.74075e-012,
  0, 0, 0, 0,
  7.490538e-014, 1.174233e-014, 5.42291e-012, 6.447455e-012,
  0, 0, 0, 0,
  1.189464e-015, 1.691791e-015, 4.122432e-012, 6.136789e-012,
  0, 0, 0, 0,
  1.31555e-015, 1.341017e-015, 4.990985e-012, 6.382807e-012,
  0, 0, 0, 0,
  1.271443e-014, 4.243659e-014, 3.072032e-012, 6.841772e-012,
  0, 0, 0, 0,
  7.48067e-014, 1.314652e-014, 6.372753e-012, 9.332739e-012,
  0, 0, 0, 0,
  8.844047e-015, 2.287604e-015, 4.130612e-012, 7.923235e-012,
  0, 0, 0, 0,
  3.849511e-014, 6.264113e-015, 4.78792e-012, 8.970056e-012,
  0, 0, 0, 0,
  5.372832e-015, 1.687487e-015, 5.938191e-012, 9.231954e-012,
  0, 0, 0, 0,
  1.298177e-015, 1.549089e-015, 3.52457e-012, 5.110972e-012,
  0, 0, 0, 0,
  2.781187e-015, 1.924865e-015, 6.282078e-012, 1.106924e-011,
  0, 0, 0, 0,
  7.086131e-015, 2.2009e-015, 1.019981e-011, 1.402387e-011,
  0, 0, 0, 0,
  1.735883e-015, 1.765689e-015, 2.646003e-012, 5.732859e-012,
  0, 0, 0, 0,
  3.095267e-015, 3.842596e-015, 5.868699e-012, 5.437831e-012,
  0, 0, 0, 0,
  3.646996e-015, 4.012981e-015, 4.391081e-012, 4.1281e-012,
  0, 0, 0, 0,
  2.424555e-015, 2.568633e-015, 6.824915e-012, 8.424729e-012,
  0, 0, 0, 0,
  2.452587e-015, 2.717092e-015, 5.09213e-012, 5.341694e-012,
  0, 0, 0, 0,
  8.749632e-015, 2.661385e-015, 5.583263e-012, 8.128617e-012,
  0, 0, 0, 0,
  1.015504e-013, 1.579873e-014, 7.385628e-012, 1.063885e-011,
  0, 0, 0, 0,
  2.156343e-015, 6.939993e-015, 7.363028e-012, 1.227591e-011,
  0, 0, 0, 0,
  1.574253e-015, 4.056339e-015, 3.803573e-012, 6.836182e-012,
  0, 0, 0, 0,
  2.646161e-015, 3.96647e-015, 5.726663e-012, 1.096652e-011,
  0, 0, 0, 0,
  8.414061e-014, 1.307427e-014, 8.319539e-012, 1.082832e-011,
  0, 0, 0, 0,
  4.740476e-015, 2.365026e-015, 8.684432e-012, 1.028301e-011,
  0, 0, 0, 0,
  3.26328e-015, 4.350498e-015, 9.703035e-012, 1.060962e-011,
  0, 0, 0, 0,
  1.092042e-015, 1.463079e-015, 2.942954e-012, 3.963798e-012,
  0, 0, 0, 0,
  1.685614e-015, 1.410831e-015, 1.067176e-011, 5.968876e-011,
  0, 0, 0, 0,
  2.476949e-015, 2.202891e-015, 9.184964e-012, 8.856861e-012,
  0, 0, 0, 0,
  5.747809e-015, 2.138806e-015, 5.399263e-012, 8.332186e-012,
  0, 0, 0, 0,
  3.454741e-015, 3.416373e-015, 7.840979e-012, 1.248667e-011,
  0, 0, 0, 0,
  1.402067e-014, 3.924916e-015, 8.840591e-012, 1.129011e-011,
  0, 0, 0, 0,
  1.85543e-014, 3.330375e-015, 5.657494e-012, 6.430588e-012,
  0, 0, 0, 0,
  1.965472e-015, 2.144111e-015, 4.444739e-012, 7.379629e-012,
  0, 0, 0, 0,
  8.4303e-015, 2.135563e-015, 2.717414e-012, 2.963395e-012,
  0, 0, 0, 0,
  1.297605e-014, 3.355237e-015, 4.677366e-012, 5.510398e-012,
  0, 0, 0, 0,
  6.518372e-014, 1.06903e-014, 3.859886e-012, 8.14191e-012,
  0, 0, 0, 0,
  3.218555e-015, 2.546623e-015, 5.210498e-012, 7.329562e-012,
  0, 0, 0, 0,
  1.570906e-015, 2.076043e-015, 4.473427e-012, 5.991399e-012,
  0, 0, 0, 0,
  1.898028e-015, 2.340662e-015, 4.098449e-012, 6.447624e-012,
  0, 0, 0, 0,
  8.149891e-014, 1.258977e-014, 1.824752e-012, 2.874233e-012,
  0, 0, 0, 0,
  2.713524e-015, 2.350304e-015, 8.558414e-012, 9.749507e-012,
  0, 0, 0, 0,
  1.3382e-015, 2.066163e-015, 7.71727e-012, 8.733087e-012,
  0, 0, 0, 0,
  2.098792e-015, 3.375384e-015, 5.19569e-012, 9.589189e-012,
  0, 0, 0, 0,
  2.538866e-014, 2.962576e-014, 1.272321e-011, 1.964637e-011,
  0, 0, 0, 0,
  3.989116e-015, 3.347635e-015, 1.019176e-011, 1.172804e-011,
  0, 0, 0, 0,
  4.308808e-015, 4.148954e-015, 6.50129e-012, 9.830543e-012,
  0, 0, 0, 0,
  2.206505e-015, 2.968558e-015, 6.540696e-012, 9.510898e-012,
  0, 0, 0, 0,
  4.30707e-014, 7.894522e-015, 7.308696e-012, 1.111301e-011,
  0, 0, 0, 0,
  3.24389e-014, 6.776009e-015, 8.221897e-012, 8.629417e-012,
  0, 0, 0, 0,
  2.491165e-015, 1.565292e-015, 3.28031e-012, 4.191139e-012,
  0, 0, 0, 0,
  2.126676e-015, 1.547435e-015, 5.013935e-012, 6.731966e-012,
  0, 0, 0, 0,
  2.356342e-014, 3.991152e-015, 4.428496e-012, 7.611571e-012,
  0, 0, 0, 0,
  5.900566e-014, 9.177033e-015, 9.669031e-012, 1.590982e-011,
  0, 0, 0, 0,
  1.728395e-015, 2.259383e-015, 7.798651e-012, 1.180417e-011,
  0, 0, 0, 0,
  1.10589e-015, 1.508733e-015, 2.341106e-012, 2.365732e-012,
  0, 0, 0, 0,
  1.059171e-015, 2.385356e-015, 3.545261e-012, 4.275462e-012,
  0, 0, 0, 0,
  1.486844e-015, 1.573586e-015, 3.004904e-012, 5.299914e-012,
  0, 0, 0, 0,
  1.737634e-015, 1.681534e-015, 3.793633e-012, 6.28329e-012,
  0, 0, 0, 0,
  9.681802e-016, 1.335972e-015, 5.658816e-012, 7.130313e-012,
  0, 0, 0, 0,
  1.245632e-015, 1.864888e-015, 2.73232e-012, 3.930078e-012,
  0, 0, 0, 0,
  2.493349e-014, 4.644121e-015, 5.922099e-012, 8.715867e-012,
  0, 0, 0, 0,
  1.597295e-015, 2.177055e-015, 4.952184e-012, 6.63401e-012,
  0, 0, 0, 0,
  2.624753e-015, 3.09733e-015, 5.878343e-012, 9.952745e-012,
  0, 0, 0, 0,
  5.058609e-015, 5.77026e-015, 1.419172e-011, 1.97468e-011,
  0, 0, 0, 0,
  6.022722e-014, 1.031152e-014, 5.945065e-012, 8.167931e-012,
  0, 0, 0, 0,
  1.782701e-014, 4.336894e-015, 4.890555e-012, 5.561242e-012,
  0, 0, 0, 0,
  2.479994e-015, 2.526346e-015, 1.264172e-011, 1.401656e-011,
  0, 0, 0, 0,
  1.234299e-015, 2.35603e-015, 4.269232e-012, 5.175687e-012,
  0, 0, 0, 0,
  3.287593e-014, 5.516486e-015, 4.870514e-012, 4.358134e-012,
  0, 0, 0, 0,
  4.846798e-014, 7.575676e-015, 2.528955e-012, 4.371363e-012,
  0, 0, 0, 0,
  3.076047e-015, 1.732689e-015, 4.059366e-012, 6.562831e-012,
  0, 0, 0, 0,
  1.726594e-015, 2.195495e-015, 5.137283e-012, 7.050079e-012,
  0, 0, 0, 0,
  1.197383e-015, 1.844414e-015, 3.749323e-012, 5.357643e-012,
  0, 0, 0, 0,
  2.014622e-015, 2.647486e-015, 9.417868e-012, 1.431381e-011,
  0, 0, 0, 0,
  2.517069e-015, 2.28623e-015, 1.37523e-011, 1.40511e-011,
  0, 0, 0, 0,
  2.365307e-015, 2.433007e-015, 1.141421e-011, 1.405076e-011,
  0, 0, 0, 0,
  2.453707e-015, 2.935006e-015, 1.763465e-011, 1.655139e-011,
  0, 0, 0, 0,
  2.769507e-014, 4.993725e-015, 7.866004e-012, 7.879065e-012,
  0, 0, 0, 0,
  1.672047e-015, 2.66569e-015, 9.332356e-012, 1.372723e-011,
  0, 0, 0, 0,
  2.355967e-015, 2.095392e-015, 1.027989e-011, 1.570444e-011,
  0, 0, 0, 0,
  2.625161e-015, 1.374488e-015, 1.708592e-011, 1.820749e-011,
  0, 0, 0, 0,
  6.906514e-014, 1.076219e-014, 6.933963e-012, 7.54105e-012,
  0, 0, 0, 0,
  9.333536e-015, 1.640201e-015, 1.28525e-011, 1.370077e-011,
  0, 0, 0, 0,
  1.874023e-015, 1.902113e-015, 4.837524e-012, 7.397659e-012,
  0, 0, 0, 0,
  3.343706e-015, 2.777306e-015, 1.117699e-011, 1.203619e-011,
  0, 0, 0, 0,
  5.090099e-014, 8.152596e-015, 8.778773e-012, 1.328366e-011,
  0, 0, 0, 0,
  3.117262e-014, 5.130089e-015, 6.718019e-012, 6.663223e-012,
  0, 0, 0, 0,
  2.350693e-015, 1.935883e-015, 9.816552e-012, 1.089824e-011,
  0, 0, 0, 0,
  3.706964e-015, 2.387245e-015, 1.508275e-011, 1.539037e-011,
  0, 0, 0, 0,
  3.793737e-015, 3.08161e-015, 6.922584e-012, 7.00039e-012,
  0, 0, 0, 0,
  2.405306e-015, 2.665056e-015, 1.1469e-011, 1.06181e-011,
  0, 0, 0, 0,
  3.375485e-015, 2.88819e-015, 1.0034e-011, 8.780867e-012,
  0, 0, 0, 0,
  2.789083e-015, 3.50131e-015, 8.901567e-012, 1.262702e-011,
  0, 0, 0, 0,
  3.788303e-015, 3.549944e-015, 1.045913e-011, 1.510012e-011,
  0, 0, 0, 0,
  3.497367e-015, 3.482036e-015, 2.935018e-012, 4.739456e-012,
  0, 0, 0, 0,
  3.383134e-015, 3.850708e-015, 3.381014e-012, 3.722036e-012,
  0, 0, 0, 0,
  3.738105e-015, 3.715837e-015, 2.806633e-012, 3.811491e-012,
  0, 0, 0, 0,
  1.491266e-014, 4.167193e-015, 5.839156e-012, 6.294162e-012,
  0, 0, 0, 0,
  7.299734e-015, 5.184279e-015, 1.776658e-011, 2.24688e-011,
  0, 0, 0, 0,
  6.354193e-015, 3.847213e-015, 2.600152e-011, 2.404408e-011,
  0, 0, 0, 0,
  8.007498e-014, 1.33305e-014, 1.829885e-011, 3.220295e-011,
  0, 0, 0, 0,
  1.065594e-014, 5.594095e-015, 5.313412e-012, 6.58274e-012,
  0, 0, 0, 0,
  1.266805e-014, 6.858353e-015, 1.147313e-011, 1.280887e-011,
  0, 0, 0, 0,
  1.309138e-014, 8.717246e-015, 1.921934e-011, 1.91511e-011,
  0, 0, 0, 0,
  1.586997e-014, 9.083283e-015, 5.653547e-012, 8.391392e-012,
  0, 0, 0, 0,
  1.825412e-014, 1.153172e-014, 1.278855e-011, 1.57674e-011,
  0, 0, 0, 0,
  2.057532e-014, 1.010323e-014, 2.982428e-012, 6.428726e-012,
  0, 0, 0, 0,
  2.73292e-014, 1.783306e-014, 5.804629e-012, 7.410292e-012,
  0, 0, 0, 0,
  3.406649e-014, 1.357438e-014, 4.679481e-012, 6.53971e-012,
  0, 0, 0, 0,
  5.599644e-014, 1.55332e-014, 6.609534e-012, 1.053158e-011,
  0, 0, 0, 0,
  1.010602e-013, 2.212689e-014, 1.125169e-011, 1.504172e-011,
  0, 0, 0, 0,
  6.148252e-014, 2.418147e-014, 4.035671e-012, 1.038339e-011,
  0, 0, 0, 0,
  1.057091e-013, 3.480967e-014, 7.852806e-012, 1.845281e-011,
  0, 0, 0, 0,
  1.331183e-013, 8.600266e-014, 7.852733e-012, 1.367993e-011,
  0, 0, 0, 0,
  1.49129e-012, 2.457158e-013, 1.289827e-011, 4.845384e-011,
  0, 0, 0, 0,
  2.037294e-013, 6.794367e-014, 9.149482e-012, 2.717959e-011,
  0, 0, 0, 0,
  2.465158e-013, 7.987923e-014, 9.824115e-012, 3.654892e-011,
  0, 0, 0, 0,
  3.672612e-013, 1.226608e-013, 1.730743e-011, 5.548714e-011,
  0, 0, 0, 0,
  6.856045e-013, 2.019201e-013, 2.557942e-011, 1.049335e-010,
  0, 0, 0, 0,
  1.176017e-012, 2.913464e-013, 1.392014e-010, 4.972024e-010,
  0, 0, 0, 0,
  1.758853e-012, 7.541959e-013, 8.456853e-011, 4.168242e-010,
  0, 0, 0, 0,
  2.565168e-012, 1.143615e-012, 1.742808e-010, 5.734656e-010,
  0, 0, 0, 0,
  4.380112e-012, 2.340361e-012, 7.782949e-010, 1.623474e-009,
  0, 0, 0, 0,
  1.265052e-011, 4.9532e-012, 1.57073e-009, 7.960697e-009,
  0, 0, 0, 0,
  1.190844e-011, 3.848853e-012, 7.948554e-010, 2.006785e-009,
  0, 0, 0, 0,
  3.739088e-012, 2.354764e-012, 6.517639e-010, 1.069036e-009,
  0, 0, 0, 0,
  1.200007e-011, 3.50951e-012, 8.7824e-010, 2.08462e-009,
  0, 0, 0, 0,
  1.339786e-011, 4.738043e-012, 8.013499e-010, 2.605253e-009,
  0, 0, 0, 0,
  3.086374e-012, 2.368344e-012, 3.491499e-010, 1.300194e-009,
  0, 0, 0, 0,
  2.538999e-012, 7.088625e-013, 1.176096e-010, 4.897829e-010,
  0, 0, 0, 0,
  1.502727e-012, 4.8114e-013, 6.093463e-011, 2.44775e-010,
  0, 0, 0, 0,
  9.876594e-013, 2.849803e-013, 3.649142e-011, 1.560628e-010,
  0, 0, 0, 0,
  5.914977e-013, 1.795224e-013, 2.48869e-011, 1.069865e-010,
  0, 0, 0, 0,
  3.698031e-013, 1.636525e-013, 2.219825e-011, 7.650081e-011,
  0, 0, 0, 0,
  2.63332e-013, 1.397212e-013, 1.671148e-011, 5.930345e-011,
  0, 0, 0, 0,
  1.947823e-013, 8.29833e-014, 1.670565e-011, 3.928647e-011,
  0, 0, 0, 0,
  1.690878e-013, 5.87818e-014, 1.406276e-011, 2.426047e-011,
  0, 0, 0, 0,
  1.138784e-013, 3.304276e-014, 1.034313e-011, 1.636237e-011,
  0, 0, 0, 0,
  7.227803e-014, 2.459901e-014, 1.056408e-011, 1.582454e-011,
  0, 0, 0, 0,
  1.116053e-013, 2.629907e-014, 8.426849e-012, 2.063596e-011,
  0, 0, 0, 0,
  5.359051e-014, 2.88836e-014, 1.526487e-011, 1.417122e-011,
  0, 0, 0, 0,
  4.725403e-014, 2.125877e-014, 6.214416e-012, 8.937994e-012,
  0, 0, 0, 0,
  2.816574e-014, 1.250196e-014, 9.22104e-012, 1.102899e-011,
  0, 0, 0, 0,
  3.057341e-014, 1.599001e-014, 1.129254e-011, 1.335523e-011,
  0, 0, 0, 0,
  3.047865e-014, 1.003243e-014, 1.281906e-011, 1.682763e-011,
  0, 0, 0, 0,
  3.09714e-014, 1.106955e-014, 1.488715e-011, 2.284411e-011,
  0, 0, 0, 0,
  2.500639e-014, 8.830091e-015, 1.989805e-011, 2.397927e-011,
  0, 0, 0, 0,
  1.637388e-014, 6.693074e-015, 1.487738e-011, 2.316287e-011,
  0, 0, 0, 0,
  6.722876e-014, 2.455479e-014, 1.803917e-011, 2.707127e-011,
  0, 0, 0, 0,
  1.481963e-014, 5.572016e-015, 1.502785e-011, 2.05502e-011,
  0, 0, 0, 0,
  8.110213e-015, 3.713652e-015, 1.861474e-011, 1.790007e-011,
  0, 0, 0, 0,
  8.132379e-015, 3.676115e-015, 1.148002e-011, 1.659701e-011,
  0, 0, 0, 0,
  6.258708e-015, 4.061571e-015, 1.504501e-011, 1.736845e-011,
  0, 0, 0, 0,
  8.080875e-015, 6.985752e-015, 1.241484e-011, 1.564691e-011,
  0, 0, 0, 0,
  6.413509e-015, 3.999656e-015, 1.566097e-011, 1.618054e-011,
  0, 0, 0, 0,
  5.300578e-015, 4.011195e-015, 9.429192e-012, 1.134126e-011,
  0, 0, 0, 0,
  2.676141e-015, 3.977793e-015, 7.391561e-012, 1.135411e-011,
  0, 0, 0, 0,
  3.631306e-015, 2.826698e-015, 7.115704e-012, 8.908319e-012,
  0, 0, 0, 0,
  4.082311e-015, 1.441141e-015, 8.725348e-012, 1.083976e-011,
  0, 0, 0, 0,
  2.691332e-015, 2.963506e-015, 6.526416e-012, 9.01678e-012,
  0, 0, 0, 0,
  2.042314e-015, 2.711773e-015, 6.831557e-012, 9.864775e-012,
  0, 0, 0, 0,
  1.812347e-015, 2.22551e-015, 6.34407e-012, 8.004733e-012,
  0, 0, 0, 0,
  2.122402e-015, 2.516501e-015, 1.075717e-011, 1.588975e-011,
  0, 0, 0, 0,
  3.020056e-015, 2.154362e-015, 1.420613e-011, 1.960583e-011,
  0, 0, 0, 0,
  2.998569e-015, 5.849917e-015, 1.839164e-011, 3.678931e-011,
  0, 0, 0, 0,
  2.72311e-014, 5.894278e-015, 2.192701e-011, 2.865685e-011,
  0, 0, 0, 0,
  2.341869e-015, 7.172523e-015, 2.00804e-011, 3.039775e-011,
  0, 0, 0, 0,
  2.579588e-015, 4.775206e-015, 1.669005e-011, 2.341632e-011,
  0, 0, 0, 0,
  2.837185e-015, 2.164503e-015, 1.014522e-011, 1.317703e-011,
  0, 0, 0, 0,
  6.334243e-014, 1.001167e-014, 7.739582e-012, 1.152237e-011,
  0, 0, 0, 0,
  1.037282e-014, 2.258948e-015, 8.628049e-012, 1.488099e-011,
  0, 0, 0, 0,
  1.667353e-015, 1.990419e-015, 9.853203e-012, 1.265135e-011,
  0, 0, 0, 0,
  1.488831e-015, 1.823764e-015, 1.19563e-011, 1.326244e-011,
  0, 0, 0, 0,
  4.661844e-014, 7.527687e-015, 1.634299e-011, 1.766711e-011,
  0, 0, 0, 0,
  3.058096e-014, 5.219302e-015, 6.859732e-012, 1.021565e-011,
  0, 0, 0, 0,
  6.252399e-015, 2.616906e-015, 1.836514e-011, 1.96303e-011,
  0, 0, 0, 0,
  2.577465e-015, 2.741487e-015, 1.556813e-011, 1.618848e-011,
  0, 0, 0, 0,
  5.86366e-015, 3.379332e-015, 1.792177e-011, 2.3388e-011,
  0, 0, 0, 0,
  2.603381e-015, 2.41146e-015, 1.983451e-011, 2.558851e-011,
  0, 0, 0, 0,
  3.083695e-015, 5.980602e-015, 2.118592e-011, 2.174609e-011,
  0, 0, 0, 0,
  3.064534e-015, 2.284496e-015, 1.309671e-011, 2.164639e-011,
  0, 0, 0, 0,
  3.04882e-015, 3.697018e-015, 1.805101e-011, 2.379967e-011,
  0, 0, 0, 0,
  2.631177e-014, 4.899504e-015, 1.834131e-011, 2.220885e-011,
  0, 0, 0, 0,
  3.080686e-015, 2.916619e-015, 2.853166e-011, 3.749712e-011,
  0, 0, 0, 0,
  3.23306e-015, 2.396597e-015, 1.646577e-011, 2.298621e-011,
  0, 0, 0, 0,
  1.717327e-015, 3.10755e-015, 1.370705e-011, 1.651363e-011,
  0, 0, 0, 0,
  6.848684e-014, 1.066425e-014, 1.028524e-011, 1.31375e-011,
  0, 0, 0, 0,
  4.083143e-015, 1.772534e-015, 6.49997e-012, 1.076787e-011,
  0, 0, 0, 0,
  2.293689e-015, 1.681595e-015, 1.367806e-011, 1.620285e-011,
  0, 0, 0, 0,
  2.366601e-015, 1.590851e-015, 1.421554e-011, 1.772278e-011,
  0, 0, 0, 0,
  5.741664e-014, 8.955707e-015, 7.478072e-012, 7.986264e-012,
  0, 0, 0, 0,
  1.96296e-014, 3.240008e-015, 1.064196e-011, 1.343874e-011,
  0, 0, 0, 0,
  1.683217e-015, 1.772863e-015, 7.472117e-012, 1.079541e-011,
  0, 0, 0, 0,
  1.456115e-015, 1.481441e-015, 5.433533e-012, 6.43125e-012,
  0, 0, 0, 0,
  1.857754e-015, 1.508157e-015, 1.104532e-011, 1.190489e-011,
  0, 0, 0, 0,
  2.014725e-015, 1.400362e-015, 7.584629e-012, 1.100456e-011,
  0, 0, 0, 0,
  1.279532e-015, 1.627681e-015, 7.788879e-012, 1.292533e-011,
  0, 0, 0, 0,
  1.479155e-015, 1.579037e-015, 1.046871e-011, 1.426415e-011,
  0, 0, 0, 0,
  4.85647e-015, 2.012845e-015, 1.19464e-011, 1.514438e-011,
  0, 0, 0, 0,
  2.559772e-014, 4.314078e-015, 1.137209e-011, 1.253991e-011,
  0, 0, 0, 0,
  1.755623e-015, 1.98237e-015, 1.662942e-011, 1.662061e-011,
  0, 0, 0, 0,
  2.210987e-015, 6.083756e-015, 1.552878e-011, 2.575001e-011,
  0, 0, 0, 0,
  2.058499e-015, 3.717979e-015, 2.150063e-011, 2.975365e-011,
  0, 0, 0, 0,
  7.267629e-014, 1.173311e-014, 2.014304e-011, 2.608495e-011,
  0, 0, 0, 0,
  4.280319e-015, 3.828978e-015, 1.904677e-011, 3.067055e-011,
  0, 0, 0, 0,
  3.188802e-015, 9.802206e-015, 4.309023e-011, 6.120407e-011,
  0, 0, 0, 0,
  4.531586e-015, 4.111708e-015, 2.262826e-011, 3.165537e-011,
  0, 0, 0, 0,
  6.712058e-014, 1.092906e-014, 2.188272e-011, 4.208102e-011,
  0, 0, 0, 0,
  1.347016e-014, 3.249652e-015, 1.692441e-011, 2.348311e-011,
  0, 0, 0, 0,
  3.474111e-015, 3.096111e-015, 2.339562e-011, 3.961852e-011,
  0, 0, 0, 0,
  3.232892e-015, 2.993939e-015, 2.066906e-011, 2.387106e-011,
  0, 0, 0, 0,
  1.689441e-014, 3.818527e-015, 3.166073e-011, 4.162662e-011,
  0, 0, 0, 0,
  1.362621e-014, 3.183952e-015, 2.070716e-011, 3.288579e-011,
  0, 0, 0, 0,
  3.492965e-015, 4.426859e-015, 3.008649e-011, 4.765159e-011,
  0, 0, 0, 0,
  2.632077e-015, 4.751394e-015, 2.40953e-011, 3.585906e-011,
  0, 0, 0, 0,
  2.302116e-014, 4.554751e-015, 2.6553e-011, 3.923646e-011,
  0, 0, 0, 0,
  5.318446e-014, 8.403018e-015, 2.295374e-011, 2.983087e-011,
  0, 0, 0, 0,
  2.214234e-015, 2.878395e-015, 1.309141e-011, 2.712574e-011,
  0, 0, 0, 0,
  1.80371e-015, 1.79359e-015, 1.311843e-011, 1.72378e-011,
  0, 0, 0, 0,
  3.114095e-015, 2.082896e-015, 1.182965e-011, 1.244159e-011,
  0, 0, 0, 0,
  7.348652e-014, 1.147986e-014, 1.837347e-011, 2.257718e-011,
  0, 0, 0, 0,
  1.360933e-015, 1.867075e-015, 1.552508e-011, 2.083357e-011,
  0, 0, 0, 0,
  1.406978e-015, 1.481064e-015, 8.137517e-012, 1.2914e-011,
  0, 0, 0, 0,
  1.695944e-015, 1.402159e-015, 9.722477e-012, 1.104292e-011,
  0, 0, 0, 0,
  1.840508e-015, 2.125488e-015, 8.140814e-012, 8.905376e-012,
  0, 0, 0, 0,
  1.520177e-015, 2.282335e-015, 1.053121e-011, 1.255778e-011,
  0, 0, 0, 0,
  1.721879e-015, 3.179505e-015, 5.389791e-012, 6.068868e-012,
  0, 0, 0, 0,
  2.110441e-014, 3.988525e-015, 1.090562e-011, 1.291366e-011,
  0, 0, 0, 0,
  5.087138e-014, 7.90284e-015, 1.231557e-011, 1.192997e-011,
  0, 0, 0, 0,
  2.417979e-014, 4.059399e-015, 1.13282e-011, 1.773344e-011,
  0, 0, 0, 0,
  8.028157e-014, 1.248114e-014, 1.196595e-011, 1.382708e-011,
  0, 0, 0, 0,
  1.700299e-014, 3.156143e-015, 1.259021e-011, 1.600274e-011,
  0, 0, 0, 0,
  2.687121e-014, 4.285376e-015, 7.941686e-012, 1.124167e-011,
  0, 0, 0, 0,
  5.284016e-014, 8.288029e-015, 1.023014e-011, 1.448015e-011,
  0, 0, 0, 0,
  2.701565e-015, 2.35227e-015, 1.052259e-011, 1.678057e-011,
  0, 0, 0, 0,
  3.181821e-015, 1.950064e-015, 8.750229e-012, 1.295271e-011,
  0, 0, 0, 0,
  2.620865e-015, 1.993323e-015, 9.726527e-012, 1.388486e-011,
  0, 0, 0, 0,
  2.542452e-015, 1.957542e-015, 1.642197e-011, 2.226014e-011,
  0, 0, 0, 0,
  1.837909e-015, 3.148045e-015, 9.654665e-012, 1.407631e-011,
  0, 0, 0, 0,
  1.554389e-015, 1.611706e-015, 1.23873e-011, 1.251248e-011,
  0, 0, 0, 0,
  2.263338e-015, 1.610117e-015, 1.863868e-011, 2.44649e-011,
  0, 0, 0, 0,
  7.192125e-014, 1.131399e-014, 1.694164e-011, 1.999655e-011,
  0, 0, 0, 0,
  3.370541e-015, 3.257157e-015, 2.211419e-011, 2.186498e-011,
  0, 0, 0, 0,
  3.359757e-015, 3.23942e-015, 2.730563e-011, 3.97049e-011,
  0, 0, 0, 0,
  3.646437e-015, 2.211057e-015, 2.367065e-011, 2.599453e-011,
  0, 0, 0, 0,
  5.975786e-014, 1.022695e-014, 3.648653e-011, 3.769442e-011,
  0, 0, 0, 0,
  2.097302e-014, 4.617023e-015, 2.415661e-011, 3.781712e-011,
  0, 0, 0, 0,
  4.056009e-015, 3.493498e-015, 2.385241e-011, 3.268037e-011,
  0, 0, 0, 0,
  3.379417e-015, 4.362558e-015, 2.334225e-011, 3.380715e-011,
  0, 0, 0, 0,
  6.71383e-015, 3.622673e-015, 4.006528e-011, 6.011164e-011,
  0, 0, 0, 0,
  2.531603e-015, 3.321215e-015, 2.880583e-011, 3.88565e-011,
  0, 0, 0, 0,
  2.321208e-015, 1.896641e-015, 1.449498e-011, 2.236828e-011,
  0, 0, 0, 0,
  2.756518e-015, 2.141078e-015, 1.760597e-011, 2.195365e-011,
  0, 0, 0, 0,
  1.242071e-014, 2.916177e-015, 1.130242e-011, 1.559055e-011,
  0, 0, 0, 0,
  6.522188e-014, 1.015064e-014, 1.109154e-011, 1.471023e-011,
  0, 0, 0, 0,
  2.337338e-015, 1.661757e-015, 1.501577e-011, 1.435712e-011,
  0, 0, 0, 0,
  1.81273e-015, 1.673469e-015, 9.693311e-012, 1.303912e-011,
  0, 0, 0, 0,
  1.663491e-015, 2.097797e-015, 1.26997e-011, 2.031546e-011,
  0, 0, 0, 0,
  7.344011e-014, 1.1398e-014, 1.280544e-011, 1.632469e-011,
  0, 0, 0, 0,
  1.605088e-015, 2.307193e-015, 1.088228e-011, 1.401075e-011,
  0, 0, 0, 0,
  2.771316e-015, 2.674617e-015, 1.549412e-011, 2.032158e-011,
  0, 0, 0, 0,
  2.642166e-015, 6.702703e-015, 1.473168e-011, 2.307607e-011,
  0, 0, 0, 0,
  2.950727e-015, 2.505622e-015, 1.279775e-011, 2.176066e-011,
  0, 0, 0, 0,
  1.589577e-015, 2.626367e-015, 2.297615e-011, 2.918971e-011,
  0, 0, 0, 0,
  2.250641e-015, 5.226189e-015, 2.6336e-011, 3.574221e-011,
  0, 0, 0, 0,
  3.857827e-015, 6.637819e-015, 2.861504e-011, 3.630543e-011,
  0, 0, 0, 0,
  3.394535e-015, 3.698712e-015, 2.404161e-011, 3.232214e-011,
  0, 0, 0, 0,
  3.340686e-015, 3.545301e-015, 1.823868e-011, 1.541947e-011,
  0, 0, 0, 0,
  2.720705e-015, 2.766824e-015, 2.037866e-011, 2.62095e-011,
  0, 0, 0, 0,
  2.341751e-015, 6.263463e-015, 1.822048e-011, 2.051245e-011,
  0, 0, 0, 0,
  1.85649e-014, 4.156846e-015, 2.453291e-011, 2.161369e-011,
  0, 0, 0, 0,
  5.685681e-014, 9.256882e-015, 1.883052e-011, 2.028171e-011,
  0, 0, 0, 0,
  2.030635e-015, 2.544589e-015, 2.319574e-011, 2.289562e-011,
  0, 0, 0, 0,
  3.00518e-015, 2.686279e-015, 1.882746e-011, 2.234363e-011,
  0, 0, 0, 0,
  5.085489e-015, 2.925181e-015, 1.798279e-011, 2.675008e-011,
  0, 0, 0, 0,
  7.397045e-014, 1.169109e-014, 1.368395e-011, 2.120577e-011,
  0, 0, 0, 0,
  2.866585e-015, 3.357791e-015, 1.155531e-011, 1.270764e-011,
  0, 0, 0, 0,
  1.45077e-015, 2.460297e-015, 1.138816e-011, 1.140979e-011,
  0, 0, 0, 0,
  1.95253e-015, 3.378812e-015, 2.410066e-011, 2.734328e-011,
  0, 0, 0, 0,
  2.263485e-015, 2.859083e-015, 1.871028e-011, 2.455118e-011,
  0, 0, 0, 0,
  1.836041e-015, 2.467524e-015, 1.92588e-011, 1.920941e-011,
  0, 0, 0, 0,
  1.400405e-015, 2.295547e-015, 1.320631e-011, 1.563093e-011,
  0, 0, 0, 0,
  2.858098e-015, 2.734211e-015, 1.471027e-011, 1.808432e-011,
  0, 0, 0, 0,
  5.716504e-014, 9.150391e-015, 1.52698e-011, 2.179155e-011,
  0, 0, 0, 0,
  1.712146e-014, 4.174344e-015, 1.56008e-011, 1.823577e-011,
  0, 0, 0, 0,
  4.162334e-015, 4.031707e-015, 2.973393e-011, 4.249465e-011,
  0, 0, 0, 0,
  4.919244e-015, 3.182695e-015, 3.326114e-011, 3.272745e-011,
  0, 0, 0, 0,
  2.922102e-014, 5.948826e-015, 1.524453e-011, 2.991266e-011,
  0, 0, 0, 0,
  5.234924e-014, 8.719667e-015, 2.889189e-011, 3.16883e-011,
  0, 0, 0, 0,
  2.907422e-015, 3.76257e-015, 2.98648e-011, 2.870617e-011,
  0, 0, 0, 0,
  2.563317e-015, 4.103907e-015, 2.438284e-011, 3.217216e-011,
  0, 0, 0, 0,
  3.193359e-015, 3.416279e-015, 1.624541e-011, 2.167796e-011,
  0, 0, 0, 0,
  3.579978e-015, 2.934812e-015, 1.312931e-011, 1.923476e-011,
  0, 0, 0, 0,
  1.831502e-015, 2.174409e-015, 1.289848e-011, 1.692982e-011,
  0, 0, 0, 0,
  2.654328e-015, 1.672896e-015, 1.59476e-011, 2.054037e-011,
  0, 0, 0, 0,
  2.163179e-015, 2.356726e-015, 1.477315e-011, 1.549319e-011,
  0, 0, 0, 0,
  7.197309e-014, 1.126751e-014, 1.677277e-011, 2.69375e-011,
  0, 0, 0, 0,
  3.52512e-015, 2.477217e-015, 2.600398e-011, 3.312563e-011,
  0, 0, 0, 0,
  3.119154e-015, 3.275416e-015, 2.228758e-011, 3.039114e-011,
  0, 0, 0, 0,
  2.307106e-015, 2.106609e-015, 1.950671e-011, 2.420964e-011,
  0, 0, 0, 0,
  6.457666e-014, 1.021122e-014, 1.96254e-011, 1.779616e-011,
  0, 0, 0, 0,
  1.286604e-014, 2.737044e-015, 1.653309e-011, 2.005056e-011,
  0, 0, 0, 0,
  2.146026e-015, 2.403535e-015, 1.919819e-011, 1.742694e-011,
  0, 0, 0, 0,
  1.912874e-015, 2.160215e-015, 2.251626e-011, 2.513084e-011,
  0, 0, 0, 0,
  2.101901e-015, 3.449786e-015, 2.206505e-011, 1.819913e-011,
  0, 0, 0, 0,
  2.064427e-015, 3.856374e-015, 1.481297e-011, 1.596802e-011,
  0, 0, 0, 0,
  5.311523e-015, 3.574278e-015, 2.127002e-011, 2.296889e-011,
  0, 0, 0, 0,
  5.568551e-015, 5.395965e-015, 3.755146e-011, 3.953458e-011,
  0, 0, 0, 0,
  6.169672e-015, 3.935438e-015, 2.310813e-011, 3.119661e-011,
  0, 0, 0, 0,
  1.644122e-014, 5.804264e-015, 2.613163e-011, 3.274503e-011,
  0, 0, 0, 0,
  5.441997e-015, 5.097875e-015, 3.046763e-011, 3.437175e-011,
  0, 0, 0, 0,
  6.286679e-015, 4.085566e-015, 1.984001e-011, 3.185343e-011,
  0, 0, 0, 0,
  4.396823e-015, 5.244467e-015, 2.638474e-011, 4.016113e-011,
  0, 0, 0, 0,
  1.708842e-015, 1.936474e-015, 2.517221e-012, 2.995015e-012,
  0, 0, 0, 0,
  1.032723e-014, 2.072516e-015, 2.25165e-011, 1.788296e-011,
  0, 0, 0, 0,
  3.617842e-014, 5.782561e-015, 4.620018e-012, 7.63601e-012,
  0, 0, 0, 0,
  6.949338e-015, 3.38687e-015, 8.502548e-012, 1.397301e-011,
  0, 0, 0, 0,
  2.508304e-015, 3.458566e-015, 4.368125e-012, 1.015293e-011,
  0, 0, 0, 0,
  1.673032e-015, 2.681079e-015, 1.23544e-011, 1.504096e-011,
  0, 0, 0, 0,
  7.459474e-014, 1.154246e-014, 5.460999e-012, 9.031149e-012,
  0, 0, 0, 0,
  1.467314e-015, 1.642659e-015, 4.85619e-012, 7.168538e-012,
  0, 0, 0, 0,
  2.096227e-015, 1.409438e-015, 5.162561e-012, 7.685829e-012,
  0, 0, 0, 0,
  1.039304e-014, 6.122978e-014, 4.64948e-012, 5.87582e-012,
  0, 0, 0, 0,
  7.386089e-014, 1.418986e-014, 4.881239e-012, 6.551863e-012,
  0, 0, 0, 0,
  8.587881e-015, 2.069972e-015, 2.772221e-012, 3.015229e-012,
  0, 0, 0, 0,
  1.212789e-014, 2.912731e-015, 4.284213e-012, 6.49566e-012,
  0, 0, 0, 0,
  2.116413e-015, 1.254869e-015, 4.157886e-012, 6.737563e-012,
  0, 0, 0, 0,
  1.534154e-015, 1.725534e-015, 4.313058e-012, 7.758708e-012,
  0, 0, 0, 0,
  2.479308e-015, 1.356763e-015, 7.847456e-012, 1.515334e-011,
  0, 0, 0, 0,
  4.955711e-015, 1.329972e-015, 1.210536e-011, 1.643473e-011,
  0, 0, 0, 0,
  1.481675e-015, 1.552255e-015, 3.046789e-012, 5.497325e-012,
  0, 0, 0, 0,
  2.995772e-015, 3.758696e-015, 4.792497e-012, 6.690604e-012,
  0, 0, 0, 0,
  2.370788e-015, 4.626124e-015, 4.112822e-012, 5.885789e-012,
  0, 0, 0, 0,
  1.456264e-015, 1.592903e-015, 3.661442e-012, 5.119138e-012,
  0, 0, 0, 0,
  1.387156e-015, 1.891534e-015, 3.441854e-012, 5.749999e-012,
  0, 0, 0, 0,
  7.753867e-015, 1.94929e-015, 6.345743e-012, 1.060547e-011,
  0, 0, 0, 0,
  7.044671e-014, 1.129484e-014, 9.748802e-012, 1.384291e-011,
  0, 0, 0, 0,
  2.722282e-015, 1.163602e-014, 8.851225e-012, 1.300901e-011,
  0, 0, 0, 0,
  1.573708e-015, 7.35609e-015, 5.818194e-012, 8.516178e-012,
  0, 0, 0, 0,
  2.266698e-015, 7.989311e-015, 6.797362e-012, 1.055289e-011,
  0, 0, 0, 0,
  8.307995e-014, 1.291142e-014, 1.091892e-011, 1.1671e-011,
  0, 0, 0, 0,
  4.056409e-015, 3.296265e-015, 4.225717e-012, 7.318828e-012,
  0, 0, 0, 0,
  1.99861e-015, 2.505242e-015, 8.427191e-012, 1.057957e-011,
  0, 0, 0, 0,
  1.39612e-015, 1.164074e-015, 3.358599e-012, 4.623374e-012,
  0, 0, 0, 0,
  2.485983e-015, 1.65829e-015, 1.20861e-011, 6.662538e-011,
  0, 0, 0, 0,
  2.610798e-015, 1.502911e-015, 6.379081e-012, 9.415754e-012,
  0, 0, 0, 0,
  7.549047e-015, 1.771621e-015, 2.93263e-012, 4.906949e-012,
  0, 0, 0, 0,
  1.98113e-015, 3.31274e-015, 7.334132e-012, 7.440263e-012,
  0, 0, 0, 0,
  2.285285e-014, 7.778233e-015, 1.064528e-011, 1.761032e-011,
  0, 0, 0, 0,
  2.758788e-014, 4.712639e-015, 4.574341e-012, 6.96159e-012,
  0, 0, 0, 0,
  2.17006e-015, 1.457552e-015, 2.422009e-012, 2.779069e-012,
  0, 0, 0, 0,
  3.510284e-015, 1.356829e-015, 2.729595e-012, 4.00185e-012,
  0, 0, 0, 0,
  1.32848e-014, 2.612708e-015, 1.61785e-012, 2.745049e-012,
  0, 0, 0, 0,
  7.689495e-014, 1.200814e-014, 2.953353e-012, 4.460171e-012,
  0, 0, 0, 0,
  5.773584e-015, 1.925937e-015, 4.841896e-012, 8.100616e-012,
  0, 0, 0, 0,
  1.523243e-015, 1.548448e-015, 3.238896e-012, 4.536286e-012,
  0, 0, 0, 0,
  1.727909e-015, 1.762242e-015, 3.955343e-012, 5.649259e-012,
  0, 0, 0, 0,
  8.036299e-014, 1.246965e-014, 2.327428e-012, 2.915354e-012,
  0, 0, 0, 0,
  2.311993e-015, 1.865756e-015, 6.735795e-012, 8.657249e-012,
  0, 0, 0, 0,
  1.101507e-015, 2.683778e-015, 7.109005e-012, 1.580767e-011,
  0, 0, 0, 0,
  1.488476e-015, 3.298601e-015, 5.438339e-012, 1.188574e-011,
  0, 0, 0, 0,
  4.334253e-014, 2.434366e-014, 6.996524e-012, 1.259836e-011,
  0, 0, 0, 0,
  6.189494e-015, 2.787136e-015, 1.262382e-011, 1.475684e-011,
  0, 0, 0, 0,
  4.351535e-015, 3.986704e-015, 6.937026e-012, 1.460762e-011,
  0, 0, 0, 0,
  1.4343e-015, 3.001038e-015, 3.872235e-012, 8.023368e-012,
  0, 0, 0, 0,
  4.267017e-014, 7.640886e-015, 6.772153e-012, 1.310166e-011,
  0, 0, 0, 0,
  3.221342e-014, 5.913917e-015, 9.028646e-012, 1.471399e-011,
  0, 0, 0, 0,
  1.352972e-015, 1.282115e-015, 2.933356e-012, 4.073325e-012,
  0, 0, 0, 0,
  1.667946e-015, 1.631059e-015, 3.102316e-012, 4.712545e-012,
  0, 0, 0, 0,
  2.210777e-014, 3.676909e-015, 5.205465e-012, 7.521816e-012,
  0, 0, 0, 0,
  5.56186e-014, 8.704392e-015, 8.306e-012, 1.100915e-011,
  0, 0, 0, 0,
  2.020854e-015, 1.312766e-015, 5.736496e-012, 7.541689e-012,
  0, 0, 0, 0,
  1.247073e-015, 9.705933e-016, 2.16887e-012, 2.084329e-012,
  0, 0, 0, 0,
  1.662495e-015, 1.097338e-015, 2.543295e-012, 5.16032e-012,
  0, 0, 0, 0,
  1.663046e-015, 1.931275e-015, 2.515344e-012, 4.946426e-012,
  0, 0, 0, 0,
  1.583628e-015, 1.024054e-015, 2.019678e-012, 2.347499e-012,
  0, 0, 0, 0,
  1.577085e-015, 1.170254e-015, 1.917983e-012, 3.666292e-012,
  0, 0, 0, 0,
  1.365514e-015, 1.388676e-015, 1.960913e-012, 2.459554e-012,
  0, 0, 0, 0,
  4.231604e-014, 7.778088e-015, 4.990478e-012, 8.033119e-012,
  0, 0, 0, 0,
  1.572099e-015, 2.144717e-015, 5.409465e-012, 7.294811e-012,
  0, 0, 0, 0,
  1.644054e-015, 2.470602e-015, 5.189005e-012, 1.086391e-011,
  0, 0, 0, 0,
  2.014519e-015, 3.829078e-015, 1.694075e-011, 2.953687e-011,
  0, 0, 0, 0,
  5.896602e-014, 9.501314e-015, 5.446041e-012, 9.32801e-012,
  0, 0, 0, 0,
  1.729864e-014, 3.228087e-015, 4.833668e-012, 8.353951e-012,
  0, 0, 0, 0,
  1.723168e-015, 2.770068e-015, 1.131469e-011, 1.082561e-011,
  0, 0, 0, 0,
  1.903882e-015, 2.049103e-015, 4.807634e-012, 7.428196e-012,
  0, 0, 0, 0,
  3.298428e-014, 5.432112e-015, 3.266844e-012, 4.360165e-012,
  0, 0, 0, 0,
  4.84152e-014, 7.587866e-015, 2.907197e-012, 3.828029e-012,
  0, 0, 0, 0,
  1.380821e-015, 1.992284e-015, 2.508422e-012, 3.481074e-012,
  0, 0, 0, 0,
  2.683361e-015, 1.984117e-015, 4.168086e-012, 5.865692e-012,
  0, 0, 0, 0,
  2.616858e-015, 1.888511e-015, 2.485813e-012, 4.418022e-012,
  0, 0, 0, 0,
  1.892358e-015, 4.093189e-015, 7.720423e-012, 1.243695e-011,
  0, 0, 0, 0,
  1.934472e-015, 3.169178e-015, 7.453815e-012, 1.068319e-011,
  0, 0, 0, 0,
  1.060243e-015, 2.054887e-015, 7.51986e-012, 1.308731e-011,
  0, 0, 0, 0,
  2.427207e-015, 5.490276e-015, 1.404285e-011, 1.902993e-011,
  0, 0, 0, 0,
  4.607346e-014, 7.701586e-015, 7.701463e-012, 9.879737e-012,
  0, 0, 0, 0,
  1.217644e-015, 3.144224e-015, 6.402942e-012, 8.439388e-012,
  0, 0, 0, 0,
  2.394511e-015, 2.471892e-015, 1.173538e-011, 1.252236e-011,
  0, 0, 0, 0,
  1.545747e-015, 2.703481e-015, 6.155249e-012, 8.108248e-012,
  0, 0, 0, 0,
  6.782015e-014, 1.072206e-014, 5.200795e-012, 8.593701e-012,
  0, 0, 0, 0,
  9.564324e-015, 3.372707e-015, 1.051983e-011, 1.485142e-011,
  0, 0, 0, 0,
  1.587439e-015, 3.117375e-015, 6.901718e-012, 1.256711e-011,
  0, 0, 0, 0,
  2.080995e-015, 2.944913e-015, 9.042593e-012, 1.452653e-011,
  0, 0, 0, 0,
  5.07142e-014, 8.872043e-015, 5.396648e-012, 9.354725e-012,
  0, 0, 0, 0,
  3.051886e-014, 5.81173e-015, 8.888607e-012, 1.40787e-011,
  0, 0, 0, 0,
  1.331606e-015, 3.049617e-015, 8.652499e-012, 1.12027e-011,
  0, 0, 0, 0,
  3.782747e-015, 2.815589e-015, 1.848146e-011, 2.235682e-011,
  0, 0, 0, 0,
  7.379692e-015, 3.757323e-015, 5.500783e-012, 7.824032e-012,
  0, 0, 0, 0,
  1.811758e-015, 3.399025e-015, 8.750783e-012, 1.30283e-011,
  0, 0, 0, 0,
  2.530468e-015, 2.405267e-015, 5.147179e-012, 7.313363e-012,
  0, 0, 0, 0,
  2.580342e-015, 1.989897e-015, 7.129205e-012, 1.094529e-011,
  0, 0, 0, 0,
  2.360619e-015, 2.65119e-015, 5.321415e-012, 9.10226e-012,
  0, 0, 0, 0,
  2.689076e-015, 2.202094e-015, 2.051319e-012, 3.778783e-012,
  0, 0, 0, 0,
  2.686018e-015, 2.463685e-015, 2.259732e-012, 3.048089e-012,
  0, 0, 0, 0,
  3.269838e-015, 3.370984e-015, 2.108338e-012, 4.305127e-012,
  0, 0, 0, 0,
  2.431546e-014, 4.374224e-015, 7.895291e-012, 9.033847e-012,
  0, 0, 0, 0,
  6.193036e-015, 3.29863e-015, 2.465212e-011, 2.844849e-011,
  0, 0, 0, 0,
  4.442929e-015, 2.347008e-015, 2.645653e-011, 3.158556e-011,
  0, 0, 0, 0,
  8.610559e-014, 1.473556e-014, 2.259767e-011, 3.147587e-011,
  0, 0, 0, 0,
  8.198074e-015, 3.964742e-015, 5.771247e-012, 8.588766e-012,
  0, 0, 0, 0,
  1.035135e-014, 6.718043e-015, 1.264832e-011, 1.806556e-011,
  0, 0, 0, 0,
  9.393733e-015, 6.42085e-015, 1.347444e-011, 2.853492e-011,
  0, 0, 0, 0,
  2.331128e-014, 7.782044e-015, 8.090061e-012, 1.469925e-011,
  0, 0, 0, 0,
  1.968777e-014, 1.048013e-014, 6.496363e-012, 8.080796e-012,
  0, 0, 0, 0,
  2.414889e-014, 7.588607e-015, 4.835403e-012, 5.418584e-012,
  0, 0, 0, 0,
  2.846648e-014, 1.414768e-014, 5.756898e-012, 6.414071e-012,
  0, 0, 0, 0,
  3.328563e-014, 1.050072e-014, 4.026366e-012, 6.494793e-012,
  0, 0, 0, 0,
  6.935183e-014, 1.661206e-014, 5.623974e-012, 1.176306e-011,
  0, 0, 0, 0,
  6.908388e-014, 1.579923e-014, 1.44046e-011, 1.565346e-011,
  0, 0, 0, 0,
  6.379006e-014, 2.032846e-014, 5.15393e-012, 1.081299e-011,
  0, 0, 0, 0,
  8.39499e-014, 3.252159e-014, 6.126339e-012, 1.24083e-011,
  0, 0, 0, 0,
  1.565886e-013, 7.968202e-014, 5.859022e-012, 1.630359e-011,
  0, 0, 0, 0,
  1.273966e-012, 2.174515e-013, 1.253174e-011, 6.3605e-011,
  0, 0, 0, 0,
  2.172316e-013, 6.662992e-014, 9.99513e-012, 3.037931e-011,
  0, 0, 0, 0,
  3.412424e-013, 7.920137e-014, 1.051072e-011, 4.811728e-011,
  0, 0, 0, 0,
  4.263055e-013, 1.178227e-013, 1.698258e-011, 6.208464e-011,
  0, 0, 0, 0,
  7.72773e-013, 2.00036e-013, 2.739418e-011, 1.158188e-010,
  0, 0, 0, 0,
  1.214658e-012, 2.839843e-013, 1.075604e-010, 3.966115e-010,
  0, 0, 0, 0,
  1.782556e-012, 7.945362e-013, 7.334254e-011, 3.359168e-010,
  0, 0, 0, 0,
  3.00034e-012, 1.085122e-012, 1.694874e-010, 6.064078e-010,
  0, 0, 0, 0,
  4.181716e-012, 2.14424e-012, 6.580809e-010, 1.551447e-009,
  0, 0, 0, 0,
  1.295172e-011, 4.329541e-012, 1.469751e-009, 7.554032e-009,
  0, 0, 0, 0,
  1.23701e-011, 3.705651e-012, 7.580748e-010, 2.292268e-009,
  0, 0, 0, 0,
  4.319742e-012, 2.490176e-012, 5.781073e-010, 1.42794e-009,
  0, 0, 0, 0,
  1.176322e-011, 3.594746e-012, 9.569006e-010, 2.407514e-009,
  0, 0, 0, 0,
  1.283331e-011, 4.374811e-012, 8.310142e-010, 3.033632e-009,
  0, 0, 0, 0,
  3.640689e-012, 2.169734e-012, 3.375636e-010, 1.274452e-009,
  0, 0, 0, 0,
  3.15729e-012, 6.669155e-013, 1.251035e-010, 5.574161e-010,
  0, 0, 0, 0,
  1.668384e-012, 5.091834e-013, 6.220629e-011, 2.573002e-010,
  0, 0, 0, 0,
  1.141796e-012, 3.512341e-013, 4.027198e-011, 1.642834e-010,
  0, 0, 0, 0,
  8.052397e-013, 2.027351e-013, 3.079521e-011, 1.065545e-010,
  0, 0, 0, 0,
  3.915809e-013, 1.718253e-013, 1.629325e-011, 7.040032e-011,
  0, 0, 0, 0,
  2.987039e-013, 1.256777e-013, 1.412612e-011, 5.281065e-011,
  0, 0, 0, 0,
  2.2687e-013, 1.369117e-013, 1.61478e-011, 5.30269e-011,
  0, 0, 0, 0,
  1.946437e-013, 5.327901e-014, 1.221736e-011, 3.245876e-011,
  0, 0, 0, 0,
  1.425367e-013, 3.385845e-014, 1.101637e-011, 2.354215e-011,
  0, 0, 0, 0,
  1.006319e-013, 2.404234e-014, 1.169273e-011, 1.810171e-011,
  0, 0, 0, 0,
  9.024835e-014, 2.601941e-014, 9.866661e-012, 2.13381e-011,
  0, 0, 0, 0,
  6.705999e-014, 2.539177e-014, 1.044219e-011, 1.814911e-011,
  0, 0, 0, 0,
  4.868499e-014, 1.859499e-014, 1.045386e-011, 1.386495e-011,
  0, 0, 0, 0,
  3.573806e-014, 1.155149e-014, 8.883085e-012, 1.375637e-011,
  0, 0, 0, 0,
  2.720975e-014, 1.583004e-014, 1.061804e-011, 1.795918e-011,
  0, 0, 0, 0,
  3.178171e-014, 1.041888e-014, 1.13056e-011, 2.494277e-011,
  0, 0, 0, 0,
  3.095228e-014, 8.427292e-015, 1.820514e-011, 2.639428e-011,
  0, 0, 0, 0,
  2.395e-014, 8.838248e-015, 1.490786e-011, 2.617025e-011,
  0, 0, 0, 0,
  1.832033e-014, 8.283585e-015, 1.482723e-011, 1.937061e-011,
  0, 0, 0, 0,
  6.913397e-014, 1.642073e-014, 1.629516e-011, 2.806126e-011,
  0, 0, 0, 0,
  1.389733e-014, 4.934519e-015, 1.422634e-011, 1.913691e-011,
  0, 0, 0, 0,
  9.292773e-015, 3.351743e-015, 2.225104e-011, 3.14611e-011,
  0, 0, 0, 0,
  7.305622e-015, 4.560842e-015, 7.3709e-012, 1.288357e-011,
  0, 0, 0, 0,
  4.848319e-015, 5.983224e-015, 8.821884e-012, 1.333102e-011,
  0, 0, 0, 0,
  7.034659e-015, 6.67274e-015, 1.142075e-011, 1.773701e-011,
  0, 0, 0, 0,
  4.195989e-015, 4.932493e-015, 1.391258e-011, 1.722978e-011,
  0, 0, 0, 0,
  3.194797e-015, 3.975699e-015, 7.413796e-012, 1.277087e-011,
  0, 0, 0, 0,
  2.522781e-015, 5.487118e-015, 8.957695e-012, 1.071593e-011,
  0, 0, 0, 0,
  1.8762e-015, 3.294225e-015, 4.795605e-012, 8.122409e-012,
  0, 0, 0, 0,
  3.876886e-015, 3.778221e-015, 7.176751e-012, 1.07966e-011,
  0, 0, 0, 0,
  2.278968e-015, 3.997739e-015, 8.669328e-012, 1.058778e-011,
  0, 0, 0, 0,
  2.599081e-015, 2.352572e-015, 5.558878e-012, 1.055249e-011,
  0, 0, 0, 0,
  2.198035e-015, 5.382315e-015, 8.464123e-012, 9.479737e-012,
  0, 0, 0, 0,
  2.345902e-015, 5.227191e-015, 1.450389e-011, 2.139719e-011,
  0, 0, 0, 0,
  3.511472e-015, 5.104099e-015, 1.287625e-011, 2.261293e-011,
  0, 0, 0, 0,
  2.829755e-015, 5.365388e-015, 2.301306e-011, 3.376288e-011,
  0, 0, 0, 0,
  4.343399e-014, 8.845976e-015, 1.405319e-011, 2.20455e-011,
  0, 0, 0, 0,
  2.767664e-015, 1.005178e-014, 1.669379e-011, 3.111646e-011,
  0, 0, 0, 0,
  2.195897e-015, 6.391604e-015, 1.18661e-011, 1.883601e-011,
  0, 0, 0, 0,
  2.183508e-015, 5.393805e-015, 8.767933e-012, 1.246969e-011,
  0, 0, 0, 0,
  6.265167e-014, 1.109528e-014, 1.172266e-011, 2.004361e-011,
  0, 0, 0, 0,
  1.014781e-014, 4.434033e-015, 9.986543e-012, 2.208224e-011,
  0, 0, 0, 0,
  2.106568e-015, 4.279206e-015, 8.465367e-012, 1.239187e-011,
  0, 0, 0, 0,
  2.008867e-015, 5.516296e-015, 8.392912e-012, 1.356191e-011,
  0, 0, 0, 0,
  4.547867e-014, 8.812164e-015, 9.858015e-012, 1.274592e-011,
  0, 0, 0, 0,
  2.861076e-014, 6.716907e-015, 7.548103e-012, 1.206197e-011,
  0, 0, 0, 0,
  8.986574e-015, 7.759513e-015, 1.207811e-011, 1.462094e-011,
  0, 0, 0, 0,
  3.987834e-015, 4.165706e-015, 1.461055e-011, 1.912168e-011,
  0, 0, 0, 0,
  4.284027e-015, 6.162655e-015, 9.371269e-012, 2.0564e-011,
  0, 0, 0, 0,
  7.139747e-015, 5.955209e-015, 1.19189e-011, 1.968466e-011,
  0, 0, 0, 0,
  3.660238e-015, 6.888347e-015, 1.869675e-011, 3.781078e-011,
  0, 0, 0, 0,
  3.256019e-015, 5.285784e-015, 1.700638e-011, 2.751682e-011,
  0, 0, 0, 0,
  3.784489e-015, 4.632516e-015, 1.464118e-011, 2.45246e-011,
  0, 0, 0, 0,
  4.405774e-014, 7.818137e-015, 1.393959e-011, 1.638023e-011,
  0, 0, 0, 0,
  3.286703e-015, 5.823969e-015, 1.689512e-011, 2.18804e-011,
  0, 0, 0, 0,
  3.362101e-015, 6.506809e-015, 1.408564e-011, 2.239728e-011,
  0, 0, 0, 0,
  3.799429e-015, 9.990103e-015, 1.726705e-011, 2.019018e-011,
  0, 0, 0, 0,
  6.672191e-014, 1.085456e-014, 6.294941e-012, 9.427015e-012,
  0, 0, 0, 0,
  4.541879e-015, 3.99909e-015, 7.975706e-012, 1.359072e-011,
  0, 0, 0, 0,
  2.726196e-015, 4.601481e-015, 1.431782e-011, 2.178346e-011,
  0, 0, 0, 0,
  1.875969e-015, 4.003323e-015, 9.823715e-012, 1.673444e-011,
  0, 0, 0, 0,
  5.508756e-014, 9.398809e-015, 8.495436e-012, 1.508991e-011,
  0, 0, 0, 0,
  1.916517e-014, 4.106125e-015, 1.001139e-011, 1.476546e-011,
  0, 0, 0, 0,
  1.713393e-015, 4.475219e-015, 9.564933e-012, 1.575762e-011,
  0, 0, 0, 0,
  2.293381e-015, 3.863247e-015, 5.796146e-012, 8.122828e-012,
  0, 0, 0, 0,
  1.909417e-015, 3.5589e-015, 8.063802e-012, 1.148443e-011,
  0, 0, 0, 0,
  2.324367e-015, 3.199072e-015, 5.603726e-012, 7.959499e-012,
  0, 0, 0, 0,
  2.031909e-015, 3.774812e-015, 7.969558e-012, 1.137359e-011,
  0, 0, 0, 0,
  2.248441e-015, 3.431893e-015, 8.737784e-012, 1.027713e-011,
  0, 0, 0, 0,
  6.758455e-015, 5.769175e-015, 1.176279e-011, 1.705666e-011,
  0, 0, 0, 0,
  3.989085e-014, 8.653325e-015, 1.235568e-011, 1.848332e-011,
  0, 0, 0, 0,
  2.814211e-015, 4.308608e-015, 1.719535e-011, 2.409035e-011,
  0, 0, 0, 0,
  2.580453e-015, 1.015559e-014, 1.273379e-011, 2.227763e-011,
  0, 0, 0, 0,
  3.768101e-015, 6.275976e-015, 2.114446e-011, 2.364973e-011,
  0, 0, 0, 0,
  7.007693e-014, 1.448045e-014, 2.584946e-011, 3.542903e-011,
  0, 0, 0, 0,
  3.011912e-015, 7.523887e-015, 2.397864e-011, 3.472695e-011,
  0, 0, 0, 0,
  3.874858e-015, 1.445455e-014, 2.354485e-011, 2.543943e-011,
  0, 0, 0, 0,
  4.343901e-015, 6.654279e-015, 2.606243e-011, 3.310611e-011,
  0, 0, 0, 0,
  6.680318e-014, 1.222713e-014, 2.456522e-011, 3.296974e-011,
  0, 0, 0, 0,
  1.306231e-014, 8.973084e-015, 3.061202e-011, 4.269847e-011,
  0, 0, 0, 0,
  3.400589e-015, 6.587107e-015, 1.997229e-011, 3.433318e-011,
  0, 0, 0, 0,
  4.015784e-015, 5.793895e-015, 2.472304e-011, 3.481745e-011,
  0, 0, 0, 0,
  2.699134e-014, 7.554473e-015, 1.795256e-011, 2.774079e-011,
  0, 0, 0, 0,
  2.029924e-014, 5.304079e-015, 2.181021e-011, 3.096328e-011,
  0, 0, 0, 0,
  4.945653e-015, 9.556434e-015, 2.453243e-011, 3.378898e-011,
  0, 0, 0, 0,
  4.371026e-015, 6.587081e-015, 1.718886e-011, 1.922358e-011,
  0, 0, 0, 0,
  2.279785e-014, 5.70447e-015, 2.010287e-011, 3.183945e-011,
  0, 0, 0, 0,
  5.327635e-014, 9.883211e-015, 1.869543e-011, 2.618824e-011,
  0, 0, 0, 0,
  2.782834e-015, 5.998079e-015, 2.042274e-011, 2.79049e-011,
  0, 0, 0, 0,
  2.431869e-015, 4.286964e-015, 1.526871e-011, 2.241006e-011,
  0, 0, 0, 0,
  4.02235e-015, 4.22812e-015, 1.781956e-011, 2.847781e-011,
  0, 0, 0, 0,
  7.103793e-014, 1.170872e-014, 1.696434e-011, 2.234913e-011,
  0, 0, 0, 0,
  2.851718e-015, 3.652905e-015, 1.154098e-011, 1.527403e-011,
  0, 0, 0, 0,
  2.034353e-015, 2.40637e-015, 8.68953e-012, 1.586594e-011,
  0, 0, 0, 0,
  2.061225e-015, 3.50957e-015, 7.174207e-012, 9.427643e-012,
  0, 0, 0, 0,
  3.040815e-015, 3.747652e-015, 9.268482e-012, 1.059042e-011,
  0, 0, 0, 0,
  2.314914e-015, 3.631598e-015, 1.092077e-011, 1.485311e-011,
  0, 0, 0, 0,
  2.347289e-015, 4.311669e-015, 1.19113e-011, 1.691509e-011,
  0, 0, 0, 0,
  2.847871e-014, 5.92564e-015, 1.013462e-011, 1.466168e-011,
  0, 0, 0, 0,
  4.834558e-014, 8.307873e-015, 1.113143e-011, 1.291996e-011,
  0, 0, 0, 0,
  2.294636e-014, 6.148424e-015, 1.066364e-011, 1.441734e-011,
  0, 0, 0, 0,
  6.20502e-014, 1.126805e-014, 1.5738e-011, 2.346972e-011,
  0, 0, 0, 0,
  1.261401e-014, 4.540406e-015, 1.187041e-011, 1.729031e-011,
  0, 0, 0, 0,
  2.624896e-014, 6.055476e-015, 1.304571e-011, 1.896122e-011,
  0, 0, 0, 0,
  5.19824e-014, 8.634334e-015, 1.517371e-011, 2.224609e-011,
  0, 0, 0, 0,
  2.70802e-015, 5.732733e-015, 2.594436e-011, 3.626769e-011,
  0, 0, 0, 0,
  3.151684e-015, 4.398776e-015, 1.872528e-011, 2.567088e-011,
  0, 0, 0, 0,
  2.405983e-015, 4.762801e-015, 1.393432e-011, 2.393814e-011,
  0, 0, 0, 0,
  4.407004e-015, 6.765746e-015, 1.999391e-011, 2.473061e-011,
  0, 0, 0, 0,
  2.598141e-015, 4.05703e-015, 1.355351e-011, 1.981177e-011,
  0, 0, 0, 0,
  2.834788e-015, 3.162543e-015, 1.752521e-011, 2.786694e-011,
  0, 0, 0, 0,
  4.087662e-015, 4.353734e-015, 1.181309e-011, 1.779065e-011,
  0, 0, 0, 0,
  7.415959e-014, 1.248892e-014, 2.627235e-011, 3.094036e-011,
  0, 0, 0, 0,
  3.230249e-015, 4.165687e-015, 2.248116e-011, 3.036825e-011,
  0, 0, 0, 0,
  4.440679e-015, 6.69974e-015, 1.617701e-011, 3.133273e-011,
  0, 0, 0, 0,
  4.141173e-015, 8.556711e-015, 1.731053e-011, 2.683682e-011,
  0, 0, 0, 0,
  5.91626e-014, 1.237025e-014, 2.236762e-011, 3.518819e-011,
  0, 0, 0, 0,
  1.983194e-014, 7.081192e-015, 2.823975e-011, 3.407886e-011,
  0, 0, 0, 0,
  7.80315e-015, 6.243026e-015, 2.986356e-011, 2.74072e-011,
  0, 0, 0, 0,
  4.225882e-015, 1.046513e-014, 2.295966e-011, 3.335625e-011,
  0, 0, 0, 0,
  6.09988e-015, 9.204704e-015, 3.401772e-011, 6.284844e-011,
  0, 0, 0, 0,
  5.183711e-015, 5.852323e-015, 2.847847e-011, 3.568616e-011,
  0, 0, 0, 0,
  4.360975e-015, 5.09689e-015, 1.890611e-011, 2.771768e-011,
  0, 0, 0, 0,
  2.554995e-015, 5.942086e-015, 1.959468e-011, 2.603267e-011,
  0, 0, 0, 0,
  1.201588e-014, 5.984708e-015, 1.519132e-011, 1.964256e-011,
  0, 0, 0, 0,
  6.350523e-014, 1.029313e-014, 1.897333e-011, 2.400329e-011,
  0, 0, 0, 0,
  2.511342e-015, 3.548402e-015, 1.101295e-011, 1.572296e-011,
  0, 0, 0, 0,
  3.39465e-015, 4.269592e-015, 1.361218e-011, 1.874628e-011,
  0, 0, 0, 0,
  2.991859e-015, 4.507582e-015, 1.756772e-011, 2.308965e-011,
  0, 0, 0, 0,
  7.208233e-014, 1.187969e-014, 1.632378e-011, 2.373285e-011,
  0, 0, 0, 0,
  3.076597e-015, 3.370043e-015, 1.47741e-011, 1.900387e-011,
  0, 0, 0, 0,
  4.15774e-015, 4.224094e-015, 1.433704e-011, 2.095138e-011,
  0, 0, 0, 0,
  4.700513e-015, 8.338095e-015, 2.665806e-011, 3.585439e-011,
  0, 0, 0, 0,
  3.169659e-015, 4.78262e-015, 2.212433e-011, 2.726049e-011,
  0, 0, 0, 0,
  3.25296e-015, 3.617195e-015, 1.571853e-011, 2.120659e-011,
  0, 0, 0, 0,
  3.303099e-015, 6.516016e-015, 1.992471e-011, 2.566401e-011,
  0, 0, 0, 0,
  5.065977e-015, 7.656425e-015, 2.170292e-011, 2.574456e-011,
  0, 0, 0, 0,
  3.813483e-015, 4.508623e-015, 1.713252e-011, 2.493889e-011,
  0, 0, 0, 0,
  5.101746e-015, 5.544235e-015, 2.41225e-011, 3.02737e-011,
  0, 0, 0, 0,
  3.752224e-015, 4.821536e-015, 1.531013e-011, 1.929392e-011,
  0, 0, 0, 0,
  4.558959e-015, 8.3861e-015, 1.915251e-011, 2.719707e-011,
  0, 0, 0, 0,
  1.842224e-014, 8.855112e-015, 2.055451e-011, 2.403095e-011,
  0, 0, 0, 0,
  5.501056e-014, 1.026177e-014, 2.717681e-011, 3.353307e-011,
  0, 0, 0, 0,
  2.613241e-015, 7.155454e-015, 2.436452e-011, 3.594527e-011,
  0, 0, 0, 0,
  2.876148e-015, 6.778349e-015, 1.651587e-011, 3.060461e-011,
  0, 0, 0, 0,
  4.844771e-015, 5.854551e-015, 2.609932e-011, 3.323068e-011,
  0, 0, 0, 0,
  7.225183e-014, 1.19927e-014, 1.967563e-011, 2.715741e-011,
  0, 0, 0, 0,
  2.455142e-015, 6.670907e-015, 1.870077e-011, 2.775615e-011,
  0, 0, 0, 0,
  2.904878e-015, 6.304105e-015, 1.993109e-011, 2.842811e-011,
  0, 0, 0, 0,
  3.382389e-015, 7.013501e-015, 2.074608e-011, 2.910494e-011,
  0, 0, 0, 0,
  5.129668e-015, 6.999901e-015, 1.854324e-011, 2.197974e-011,
  0, 0, 0, 0,
  2.947853e-015, 6.065917e-015, 2.048517e-011, 2.645085e-011,
  0, 0, 0, 0,
  2.237586e-015, 6.126918e-015, 1.704884e-011, 2.314607e-011,
  0, 0, 0, 0,
  3.201556e-015, 5.21156e-015, 2.13712e-011, 2.926067e-011,
  0, 0, 0, 0,
  5.80071e-014, 1.049631e-014, 1.392127e-011, 2.653755e-011,
  0, 0, 0, 0,
  1.788262e-014, 6.998533e-015, 1.934893e-011, 2.858841e-011,
  0, 0, 0, 0,
  6.496963e-015, 6.114676e-015, 3.049324e-011, 3.688578e-011,
  0, 0, 0, 0,
  6.160262e-015, 6.261505e-015, 3.059e-011, 4.393218e-011,
  0, 0, 0, 0,
  2.859598e-014, 7.285341e-015, 2.543357e-011, 3.167807e-011,
  0, 0, 0, 0,
  5.290003e-014, 1.195862e-014, 3.179986e-011, 4.10819e-011,
  0, 0, 0, 0,
  5.894404e-015, 7.864522e-015, 1.61934e-011, 2.042345e-011,
  0, 0, 0, 0,
  8.239655e-015, 1.183095e-014, 3.215469e-011, 4.284133e-011,
  0, 0, 0, 0,
  4.422553e-015, 9.543525e-015, 2.568886e-011, 3.055754e-011,
  0, 0, 0, 0,
  4.875673e-015, 5.115339e-015, 1.357764e-011, 1.810383e-011,
  0, 0, 0, 0,
  3.321548e-015, 4.818365e-015, 2.381243e-011, 3.315343e-011,
  0, 0, 0, 0,
  2.069264e-015, 5.453573e-015, 1.86529e-011, 2.82328e-011,
  0, 0, 0, 0,
  3.523183e-015, 6.830035e-015, 2.84287e-011, 3.561089e-011,
  0, 0, 0, 0,
  7.057599e-014, 1.245839e-014, 1.87191e-011, 2.927211e-011,
  0, 0, 0, 0,
  3.050229e-015, 6.106333e-015, 1.940845e-011, 2.12417e-011,
  0, 0, 0, 0,
  3.781352e-015, 5.600556e-015, 1.859457e-011, 2.129012e-011,
  0, 0, 0, 0,
  2.925033e-015, 7.136304e-015, 2.171196e-011, 2.238257e-011,
  0, 0, 0, 0,
  6.314772e-014, 1.142095e-014, 2.958974e-011, 3.884612e-011,
  0, 0, 0, 0,
  1.290217e-014, 5.527936e-015, 1.780573e-011, 2.364911e-011,
  0, 0, 0, 0,
  4.090322e-015, 8.444199e-015, 1.589278e-011, 3.056862e-011,
  0, 0, 0, 0,
  4.470775e-015, 4.382198e-015, 2.522966e-011, 3.549702e-011,
  0, 0, 0, 0,
  4.646098e-015, 5.213214e-015, 1.749786e-011, 2.2229e-011,
  0, 0, 0, 0,
  3.850985e-015, 7.225942e-015, 2.962689e-011, 2.908184e-011,
  0, 0, 0, 0,
  5.367312e-015, 6.098795e-015, 2.054529e-011, 2.028849e-011,
  0, 0, 0, 0,
  6.036015e-015, 6.551032e-015, 3.808963e-011, 4.161855e-011,
  0, 0, 0, 0,
  1.047787e-014, 5.404629e-015, 2.204601e-011, 3.677703e-011,
  0, 0, 0, 0,
  2.781217e-014, 7.323033e-015, 2.476619e-011, 3.587293e-011,
  0, 0, 0, 0,
  5.918176e-015, 8.25257e-015, 3.352809e-011, 4.037022e-011,
  0, 0, 0, 0,
  7.959086e-015, 7.726025e-015, 2.744837e-011, 3.412022e-011,
  0, 0, 0, 0,
  6.256641e-015, 6.404164e-015, 3.729291e-011, 6.156524e-011,
  0, 0, 0, 0,
  2.749599e-015, 2.018595e-015, 5.161922e-012, 4.957559e-012,
  0, 0, 0, 0,
  1.503022e-014, 3.237063e-015, 3.091406e-011, 2.596146e-011,
  0, 0, 0, 0,
  4.921347e-014, 7.874542e-015, 5.606478e-012, 5.378983e-012,
  0, 0, 0, 0,
  4.474301e-015, 4.089077e-015, 9.618494e-012, 2.356522e-011,
  0, 0, 0, 0,
  2.31755e-015, 3.190306e-015, 5.491609e-012, 8.639709e-012,
  0, 0, 0, 0,
  2.112521e-015, 2.651472e-015, 1.16198e-011, 1.91957e-011,
  0, 0, 0, 0,
  7.418596e-014, 1.164716e-014, 7.11013e-012, 8.236711e-012,
  0, 0, 0, 0,
  1.990224e-015, 2.026563e-015, 4.461811e-012, 6.397991e-012,
  0, 0, 0, 0,
  3.955503e-015, 2.4792e-015, 7.198491e-012, 5.563579e-012,
  0, 0, 0, 0,
  8.858833e-015, 5.066065e-014, 5.536085e-012, 5.157387e-012,
  0, 0, 0, 0,
  7.428113e-014, 1.378203e-014, 5.036143e-012, 7.814982e-012,
  0, 0, 0, 0,
  8.75691e-015, 1.960611e-015, 3.407429e-012, 4.728109e-012,
  0, 0, 0, 0,
  4.068931e-015, 2.289926e-015, 5.115271e-012, 4.893632e-012,
  0, 0, 0, 0,
  1.593695e-015, 1.402745e-015, 4.42241e-012, 4.876986e-012,
  0, 0, 0, 0,
  2.331531e-015, 1.767063e-015, 3.290389e-012, 5.492024e-012,
  0, 0, 0, 0,
  2.212992e-015, 1.823591e-015, 3.826551e-012, 4.837421e-012,
  0, 0, 0, 0,
  6.775926e-015, 2.295734e-015, 1.016066e-011, 1.672144e-011,
  0, 0, 0, 0,
  1.901796e-015, 1.838625e-015, 2.911203e-012, 3.998441e-012,
  0, 0, 0, 0,
  2.584375e-015, 5.637884e-015, 3.022019e-012, 5.304164e-012,
  0, 0, 0, 0,
  2.048674e-015, 2.605409e-015, 3.62381e-012, 5.924412e-012,
  0, 0, 0, 0,
  1.815722e-015, 2.164809e-015, 6.84614e-012, 8.199812e-012,
  0, 0, 0, 0,
  2.33742e-015, 1.82318e-015, 6.746608e-012, 8.348188e-012,
  0, 0, 0, 0,
  7.759744e-015, 2.268753e-015, 6.323163e-012, 7.502665e-012,
  0, 0, 0, 0,
  8.455726e-014, 1.305555e-014, 6.821798e-012, 8.220819e-012,
  0, 0, 0, 0,
  3.405906e-015, 1.667729e-014, 5.071493e-012, 7.375603e-012,
  0, 0, 0, 0,
  2.203786e-015, 9.22717e-015, 4.455109e-012, 5.080228e-012,
  0, 0, 0, 0,
  4.07337e-015, 1.448692e-014, 1.125032e-011, 1.672765e-011,
  0, 0, 0, 0,
  7.947552e-014, 1.28072e-014, 1.992366e-011, 2.137345e-011,
  0, 0, 0, 0,
  3.947059e-015, 3.447258e-015, 5.862459e-012, 9.779125e-012,
  0, 0, 0, 0,
  2.768851e-015, 2.487762e-015, 8.204177e-012, 1.137961e-011,
  0, 0, 0, 0,
  1.60422e-015, 1.464952e-015, 4.049117e-012, 4.454722e-012,
  0, 0, 0, 0,
  2.948281e-015, 1.708454e-015, 1.365309e-011, 7.029798e-011,
  0, 0, 0, 0,
  2.336677e-015, 1.682119e-015, 9.733075e-012, 1.049225e-011,
  0, 0, 0, 0,
  1.215168e-014, 2.308321e-015, 4.492173e-012, 5.098979e-012,
  0, 0, 0, 0,
  2.427507e-015, 1.974215e-015, 6.54234e-012, 8.772464e-012,
  0, 0, 0, 0,
  3.290283e-014, 5.889122e-015, 7.880213e-012, 1.017096e-011,
  0, 0, 0, 0,
  3.993278e-014, 6.343186e-015, 3.259972e-012, 4.1185e-012,
  0, 0, 0, 0,
  2.293393e-015, 1.769876e-015, 3.831252e-012, 3.993101e-012,
  0, 0, 0, 0,
  1.030439e-014, 2.439709e-015, 3.278762e-012, 3.508838e-012,
  0, 0, 0, 0,
  1.324638e-014, 3.13996e-015, 3.607326e-012, 3.223898e-012,
  0, 0, 0, 0,
  8.563101e-014, 1.334908e-014, 4.935401e-012, 4.814509e-012,
  0, 0, 0, 0,
  7.658132e-015, 1.903067e-015, 6.08162e-012, 7.654691e-012,
  0, 0, 0, 0,
  1.955205e-015, 1.652018e-015, 4.952631e-012, 5.037259e-012,
  0, 0, 0, 0,
  1.844236e-015, 1.850685e-015, 4.88862e-012, 7.51743e-012,
  0, 0, 0, 0,
  8.127292e-014, 1.253739e-014, 3.068415e-012, 3.317035e-012,
  0, 0, 0, 0,
  4.52244e-015, 3.300015e-015, 5.369335e-012, 6.713789e-012,
  0, 0, 0, 0,
  2.373885e-015, 3.253347e-015, 5.670713e-012, 9.737967e-012,
  0, 0, 0, 0,
  1.235953e-015, 3.897146e-015, 3.000637e-012, 4.755685e-012,
  0, 0, 0, 0,
  5.842906e-014, 2.295519e-014, 7.160571e-012, 7.957256e-012,
  0, 0, 0, 0,
  7.989293e-015, 3.127122e-015, 1.849815e-011, 1.910529e-011,
  0, 0, 0, 0,
  2.621212e-015, 3.122847e-015, 5.170545e-012, 8.525443e-012,
  0, 0, 0, 0,
  1.670229e-015, 3.265466e-015, 3.451449e-012, 3.882073e-012,
  0, 0, 0, 0,
  4.265449e-014, 7.80818e-015, 3.74121e-012, 3.945324e-012,
  0, 0, 0, 0,
  3.163443e-014, 6.790041e-015, 4.849709e-012, 5.156181e-012,
  0, 0, 0, 0,
  1.831277e-015, 1.684096e-015, 2.691196e-012, 3.289747e-012,
  0, 0, 0, 0,
  1.085133e-015, 1.364576e-015, 4.256161e-012, 4.844829e-012,
  0, 0, 0, 0,
  2.311779e-014, 3.792197e-015, 4.178253e-012, 5.01727e-012,
  0, 0, 0, 0,
  5.816698e-014, 9.199097e-015, 9.471132e-012, 1.373044e-011,
  0, 0, 0, 0,
  1.529016e-015, 2.226222e-015, 5.281151e-012, 7.053439e-012,
  0, 0, 0, 0,
  1.346017e-015, 1.59704e-015, 4.748966e-012, 4.787969e-012,
  0, 0, 0, 0,
  1.730734e-015, 1.744761e-015, 3.239599e-012, 3.411001e-012,
  0, 0, 0, 0,
  1.689153e-015, 2.011671e-015, 4.270827e-012, 4.095667e-012,
  0, 0, 0, 0,
  1.998032e-015, 1.533897e-015, 2.939734e-012, 3.562542e-012,
  0, 0, 0, 0,
  1.38008e-015, 1.463699e-015, 2.546092e-012, 3.289915e-012,
  0, 0, 0, 0,
  2.074701e-015, 1.64057e-015, 2.626446e-012, 2.733868e-012,
  0, 0, 0, 0,
  5.905794e-014, 1.042456e-014, 6.210824e-012, 1.00026e-011,
  0, 0, 0, 0,
  2.576377e-015, 2.787546e-015, 2.797307e-012, 4.071472e-012,
  0, 0, 0, 0,
  2.279885e-015, 4.489779e-015, 6.988956e-012, 8.082757e-012,
  0, 0, 0, 0,
  1.650388e-015, 5.311384e-015, 1.293024e-011, 2.17694e-011,
  0, 0, 0, 0,
  5.855307e-014, 9.333951e-015, 4.511145e-012, 6.455011e-012,
  0, 0, 0, 0,
  1.726295e-014, 3.19852e-015, 2.594465e-012, 3.56388e-012,
  0, 0, 0, 0,
  2.345261e-015, 2.545053e-015, 2.037424e-011, 2.308052e-011,
  0, 0, 0, 0,
  1.317502e-015, 1.515448e-015, 3.566466e-012, 3.575733e-012,
  0, 0, 0, 0,
  3.247273e-014, 5.316536e-015, 2.843931e-012, 3.123613e-012,
  0, 0, 0, 0,
  4.762377e-014, 7.500789e-015, 3.464245e-012, 3.705837e-012,
  0, 0, 0, 0,
  1.074574e-015, 2.022392e-015, 4.315825e-012, 4.493653e-012,
  0, 0, 0, 0,
  1.981832e-015, 1.197689e-015, 2.378953e-012, 2.749967e-012,
  0, 0, 0, 0,
  2.200793e-015, 2.71446e-015, 3.707353e-012, 4.125406e-012,
  0, 0, 0, 0,
  2.906988e-015, 5.14935e-015, 8.067933e-012, 1.654466e-011,
  0, 0, 0, 0,
  3.307987e-015, 4.221001e-015, 9.379758e-012, 1.384918e-011,
  0, 0, 0, 0,
  1.752565e-015, 2.29484e-015, 8.013968e-012, 1.240635e-011,
  0, 0, 0, 0,
  1.9917e-015, 5.007277e-015, 9.869257e-012, 1.345452e-011,
  0, 0, 0, 0,
  6.606736e-014, 1.152474e-014, 8.449249e-012, 1.105727e-011,
  0, 0, 0, 0,
  3.203467e-015, 6.757433e-015, 1.472961e-011, 2.016088e-011,
  0, 0, 0, 0,
  2.867829e-015, 2.284751e-015, 8.447282e-012, 1.599478e-011,
  0, 0, 0, 0,
  2.494711e-015, 4.31393e-015, 7.254258e-012, 9.866501e-012,
  0, 0, 0, 0,
  6.690229e-014, 1.114032e-014, 6.234891e-012, 8.923265e-012,
  0, 0, 0, 0,
  1.007555e-014, 3.652301e-015, 8.416665e-012, 1.295444e-011,
  0, 0, 0, 0,
  2.671946e-015, 4.166328e-015, 5.710461e-012, 6.929382e-012,
  0, 0, 0, 0,
  1.980622e-015, 8.20803e-015, 1.260621e-011, 2.455e-011,
  0, 0, 0, 0,
  5.112908e-014, 9.47779e-015, 1.427751e-011, 2.305442e-011,
  0, 0, 0, 0,
  3.090258e-014, 5.943119e-015, 1.009939e-011, 1.462427e-011,
  0, 0, 0, 0,
  2.29854e-015, 5.061916e-015, 1.10076e-011, 1.222004e-011,
  0, 0, 0, 0,
  3.775065e-015, 2.103164e-015, 2.090663e-011, 2.342258e-011,
  0, 0, 0, 0,
  7.51087e-015, 2.92242e-015, 5.160372e-012, 1.123021e-011,
  0, 0, 0, 0,
  1.813129e-015, 4.595643e-015, 6.04116e-012, 9.131794e-012,
  0, 0, 0, 0,
  2.316857e-015, 1.091804e-015, 5.265613e-012, 7.039271e-012,
  0, 0, 0, 0,
  2.468962e-015, 2.114189e-015, 6.979473e-012, 9.455503e-012,
  0, 0, 0, 0,
  2.016884e-015, 3.047108e-015, 7.788381e-012, 1.418042e-011,
  0, 0, 0, 0,
  2.488898e-015, 2.176509e-015, 3.890907e-012, 4.02481e-012,
  0, 0, 0, 0,
  2.801556e-015, 1.884957e-015, 4.212111e-012, 4.792704e-012,
  0, 0, 0, 0,
  2.643694e-015, 4.896196e-015, 3.125175e-012, 3.106512e-012,
  0, 0, 0, 0,
  2.68848e-014, 4.578908e-015, 1.00121e-011, 1.094227e-011,
  0, 0, 0, 0,
  5.680524e-015, 2.566296e-015, 3.08576e-011, 3.821785e-011,
  0, 0, 0, 0,
  7.69002e-015, 2.716417e-015, 3.175771e-011, 3.877927e-011,
  0, 0, 0, 0,
  5.432085e-014, 9.314141e-015, 3.03959e-011, 3.685012e-011,
  0, 0, 0, 0,
  7.408536e-015, 4.223639e-015, 4.566849e-012, 7.932428e-012,
  0, 0, 0, 0,
  1.051934e-014, 4.690853e-015, 9.386047e-012, 1.111852e-011,
  0, 0, 0, 0,
  1.392019e-014, 9.046503e-015, 2.761077e-011, 3.404184e-011,
  0, 0, 0, 0,
  1.861685e-014, 4.860297e-015, 7.308738e-012, 1.309057e-011,
  0, 0, 0, 0,
  1.540084e-014, 8.036009e-015, 7.693092e-012, 9.243319e-012,
  0, 0, 0, 0,
  3.121308e-014, 9.429798e-015, 4.214972e-012, 9.097473e-012,
  0, 0, 0, 0,
  2.491586e-014, 1.299324e-014, 3.956629e-012, 7.214837e-012,
  0, 0, 0, 0,
  4.018602e-014, 1.120954e-014, 3.7519e-012, 6.743759e-012,
  0, 0, 0, 0,
  6.993082e-014, 1.506416e-014, 6.587143e-012, 9.304807e-012,
  0, 0, 0, 0,
  7.947148e-014, 1.828126e-014, 2.012308e-011, 2.264067e-011,
  0, 0, 0, 0,
  6.601731e-014, 1.758822e-014, 4.671636e-012, 8.929427e-012,
  0, 0, 0, 0,
  1.198145e-013, 3.252763e-014, 5.912647e-012, 1.534707e-011,
  0, 0, 0, 0,
  1.385261e-013, 5.720696e-014, 5.384862e-012, 2.290901e-011,
  0, 0, 0, 0,
  8.921944e-013, 1.500235e-013, 1.090743e-011, 5.805963e-011,
  0, 0, 0, 0,
  2.391914e-013, 6.033682e-014, 8.878148e-012, 2.673291e-011,
  0, 0, 0, 0,
  6.109638e-013, 1.230397e-013, 1.817614e-011, 7.640372e-011,
  0, 0, 0, 0,
  5.382501e-013, 1.263192e-013, 2.107484e-011, 8.422673e-011,
  0, 0, 0, 0,
  1.203828e-012, 2.705164e-013, 4.217955e-011, 1.809053e-010,
  0, 0, 0, 0,
  1.758015e-012, 3.516843e-013, 1.19655e-010, 4.453494e-010,
  0, 0, 0, 0,
  2.001144e-012, 6.186042e-013, 8.563334e-011, 4.005967e-010,
  0, 0, 0, 0,
  3.248191e-012, 1.057052e-012, 1.677317e-010, 6.295113e-010,
  0, 0, 0, 0,
  5.626697e-012, 2.171699e-012, 6.34128e-010, 1.66821e-009,
  0, 0, 0, 0,
  1.297559e-011, 4.344925e-012, 1.434293e-009, 7.191128e-009,
  0, 0, 0, 0,
  1.333193e-011, 3.995937e-012, 9.343591e-010, 3.03337e-009,
  0, 0, 0, 0,
  5.949503e-012, 2.715316e-012, 6.847823e-010, 1.794281e-009,
  0, 0, 0, 0,
  1.255648e-011, 3.901533e-012, 1.0196e-009, 2.774802e-009,
  0, 0, 0, 0,
  1.315404e-011, 4.43688e-012, 7.989205e-010, 2.814415e-009,
  0, 0, 0, 0,
  3.974784e-012, 2.170032e-012, 3.592447e-010, 1.385817e-009,
  0, 0, 0, 0,
  3.391356e-012, 6.739959e-013, 1.459147e-010, 5.940398e-010,
  0, 0, 0, 0,
  1.806076e-012, 4.832987e-013, 6.74544e-011, 2.762031e-010,
  0, 0, 0, 0,
  1.226052e-012, 3.310874e-013, 4.238355e-011, 1.817865e-010,
  0, 0, 0, 0,
  8.046151e-013, 2.367162e-013, 3.461727e-011, 1.238658e-010,
  0, 0, 0, 0,
  4.068188e-013, 1.487713e-013, 1.915053e-011, 8.554689e-011,
  0, 0, 0, 0,
  3.118004e-013, 1.587383e-013, 1.939764e-011, 5.54667e-011,
  0, 0, 0, 0,
  3.131276e-013, 1.581222e-013, 2.034842e-011, 4.116407e-011,
  0, 0, 0, 0,
  2.506837e-013, 6.916004e-014, 1.826287e-011, 6.094348e-011,
  0, 0, 0, 0,
  2.383599e-013, 4.389502e-014, 1.217626e-011, 2.492014e-011,
  0, 0, 0, 0,
  8.310555e-014, 2.651573e-014, 1.222255e-011, 2.870921e-011,
  0, 0, 0, 0,
  1.150932e-013, 2.905414e-014, 1.011743e-011, 2.906085e-011,
  0, 0, 0, 0,
  7.426157e-014, 2.501388e-014, 1.552015e-011, 4.149453e-011,
  0, 0, 0, 0,
  4.095158e-014, 1.574279e-014, 8.090272e-012, 8.770334e-012,
  0, 0, 0, 0,
  4.502276e-014, 1.088237e-014, 1.174447e-011, 1.553057e-011,
  0, 0, 0, 0,
  2.764306e-014, 2.100121e-014, 1.248248e-011, 2.068755e-011,
  0, 0, 0, 0,
  3.387364e-014, 1.508426e-014, 1.707184e-011, 2.487215e-011,
  0, 0, 0, 0,
  2.141489e-014, 1.550426e-014, 1.642965e-011, 2.984944e-011,
  0, 0, 0, 0,
  2.229101e-014, 1.961392e-014, 3.073525e-011, 5.401775e-011,
  0, 0, 0, 0,
  1.786708e-014, 3.111975e-014, 1.775935e-011, 2.950173e-011,
  0, 0, 0, 0,
  7.223941e-014, 2.425167e-014, 1.991045e-011, 3.336044e-011,
  0, 0, 0, 0,
  1.20239e-014, 2.330305e-014, 1.930065e-011, 3.171774e-011,
  0, 0, 0, 0,
  6.5668e-015, 1.109031e-014, 2.15575e-011, 3.332216e-011,
  0, 0, 0, 0,
  5.924973e-015, 1.248644e-014, 1.444211e-011, 2.068611e-011,
  0, 0, 0, 0,
  5.416165e-015, 1.353029e-014, 8.750788e-012, 1.571284e-011,
  0, 0, 0, 0,
  5.297527e-015, 1.33065e-014, 9.436144e-012, 1.74704e-011,
  0, 0, 0, 0,
  4.905648e-015, 8.023095e-015, 1.812112e-011, 1.655791e-011,
  0, 0, 0, 0,
  2.579678e-015, 7.56402e-015, 7.907729e-012, 1.388593e-011,
  0, 0, 0, 0,
  2.817817e-015, 1.093132e-014, 1.966784e-011, 3.304342e-011,
  0, 0, 0, 0,
  3.353608e-015, 6.264875e-015, 7.744948e-012, 1.368153e-011,
  0, 0, 0, 0,
  2.463394e-015, 9.879557e-015, 6.527861e-012, 1.543633e-011,
  0, 0, 0, 0,
  2.690012e-015, 1.037774e-014, 7.750927e-012, 1.774004e-011,
  0, 0, 0, 0,
  5.587514e-015, 9.322323e-015, 9.63698e-012, 1.891678e-011,
  0, 0, 0, 0,
  2.886128e-015, 8.261394e-015, 1.382612e-011, 2.206221e-011,
  0, 0, 0, 0,
  3.820889e-015, 1.519596e-014, 1.4675e-011, 3.035437e-011,
  0, 0, 0, 0,
  5.61141e-015, 1.74476e-014, 1.537438e-011, 3.379885e-011,
  0, 0, 0, 0,
  8.019587e-015, 4.346361e-014, 2.091979e-011, 5.296475e-011,
  0, 0, 0, 0,
  6.011233e-014, 2.85033e-014, 2.943711e-011, 5.892877e-011,
  0, 0, 0, 0,
  6.84859e-015, 3.430574e-014, 2.579027e-011, 5.085746e-011,
  0, 0, 0, 0,
  5.502735e-015, 3.014053e-014, 1.519514e-011, 3.383837e-011,
  0, 0, 0, 0,
  4.021564e-015, 1.179256e-014, 2.098476e-011, 3.242864e-011,
  0, 0, 0, 0,
  6.289378e-014, 2.378071e-014, 2.182039e-011, 4.756748e-011,
  0, 0, 0, 0,
  1.058661e-014, 1.396359e-014, 1.676573e-011, 2.910398e-011,
  0, 0, 0, 0,
  3.914119e-015, 1.297212e-014, 8.99379e-012, 1.503906e-011,
  0, 0, 0, 0,
  3.703584e-015, 1.851038e-014, 1.647731e-011, 2.819443e-011,
  0, 0, 0, 0,
  4.682602e-014, 1.706304e-014, 1.313991e-011, 2.394082e-011,
  0, 0, 0, 0,
  2.977163e-014, 1.090945e-014, 1.185429e-011, 2.168012e-011,
  0, 0, 0, 0,
  9.791843e-015, 3.156768e-014, 1.423353e-011, 2.818235e-011,
  0, 0, 0, 0,
  5.641675e-015, 1.631048e-014, 2.14023e-011, 3.598409e-011,
  0, 0, 0, 0,
  7.43336e-015, 2.609179e-014, 1.215398e-011, 2.445887e-011,
  0, 0, 0, 0,
  6.328332e-015, 1.902687e-014, 2.356459e-011, 3.892349e-011,
  0, 0, 0, 0,
  8.808269e-015, 3.907622e-014, 2.784084e-011, 5.018349e-011,
  0, 0, 0, 0,
  6.319221e-015, 2.387109e-014, 1.850587e-011, 4.202115e-011,
  0, 0, 0, 0,
  7.382379e-015, 2.541483e-014, 3.018968e-011, 4.61529e-011,
  0, 0, 0, 0,
  6.028976e-014, 1.634831e-014, 2.670551e-011, 4.33791e-011,
  0, 0, 0, 0,
  7.331069e-015, 2.694971e-014, 3.786952e-011, 6.967972e-011,
  0, 0, 0, 0,
  7.028567e-015, 2.283871e-014, 2.424644e-011, 4.901352e-011,
  0, 0, 0, 0,
  6.608473e-015, 3.836125e-014, 2.369884e-011, 4.551552e-011,
  0, 0, 0, 0,
  6.924317e-014, 1.864539e-014, 9.675736e-012, 1.811078e-011,
  0, 0, 0, 0,
  6.031807e-015, 1.568958e-014, 1.099553e-011, 2.43667e-011,
  0, 0, 0, 0,
  3.921898e-015, 1.474126e-014, 1.170178e-011, 1.920543e-011,
  0, 0, 0, 0,
  3.240251e-015, 8.404193e-015, 1.915605e-011, 3.554289e-011,
  0, 0, 0, 0,
  5.803809e-014, 1.183687e-014, 9.887604e-012, 1.693744e-011,
  0, 0, 0, 0,
  1.919885e-014, 7.626929e-015, 9.304724e-012, 1.57728e-011,
  0, 0, 0, 0,
  2.683679e-015, 1.274383e-014, 9.880135e-012, 2.054182e-011,
  0, 0, 0, 0,
  2.824341e-015, 9.794289e-015, 8.210319e-012, 1.427282e-011,
  0, 0, 0, 0,
  3.453084e-015, 1.259981e-014, 9.977821e-012, 2.500529e-011,
  0, 0, 0, 0,
  2.277541e-015, 9.280893e-015, 1.021193e-011, 1.833102e-011,
  0, 0, 0, 0,
  3.303276e-015, 1.01708e-014, 8.932878e-012, 1.362864e-011,
  0, 0, 0, 0,
  3.245747e-015, 8.814193e-015, 1.736235e-011, 3.382503e-011,
  0, 0, 0, 0,
  1.112432e-014, 2.794282e-014, 2.346723e-011, 3.957431e-011,
  0, 0, 0, 0,
  5.537939e-014, 2.298924e-014, 2.072814e-011, 3.812612e-011,
  0, 0, 0, 0,
  4.878533e-015, 2.430876e-014, 1.750197e-011, 3.494185e-011,
  0, 0, 0, 0,
  6.148062e-015, 3.357503e-014, 2.658946e-011, 4.897169e-011,
  0, 0, 0, 0,
  7.851201e-015, 3.001846e-014, 4.239811e-011, 6.947799e-011,
  0, 0, 0, 0,
  7.182793e-014, 3.287264e-014, 4.619536e-011, 7.048249e-011,
  0, 0, 0, 0,
  9.56213e-015, 4.057457e-014, 4.225893e-011, 7.767738e-011,
  0, 0, 0, 0,
  1.187749e-014, 5.841614e-014, 4.927934e-011, 9.097516e-011,
  0, 0, 0, 0,
  9.782178e-015, 2.275833e-014, 4.556224e-011, 7.130205e-011,
  0, 0, 0, 0,
  6.479449e-014, 2.450654e-014, 6.061399e-011, 1.059469e-010,
  0, 0, 0, 0,
  1.30599e-014, 2.906229e-014, 3.522435e-011, 6.024806e-011,
  0, 0, 0, 0,
  6.891008e-015, 2.535179e-014, 4.28022e-011, 5.767298e-011,
  0, 0, 0, 0,
  8.881881e-015, 2.789156e-014, 3.647061e-011, 5.388274e-011,
  0, 0, 0, 0,
  3.668065e-014, 2.317333e-014, 5.541396e-011, 9.028626e-011,
  0, 0, 0, 0,
  2.945445e-014, 1.958929e-014, 3.605908e-011, 5.679698e-011,
  0, 0, 0, 0,
  1.086117e-014, 2.455044e-014, 5.467753e-011, 8.667273e-011,
  0, 0, 0, 0,
  7.489935e-015, 2.810029e-014, 5.722644e-011, 1.027838e-010,
  0, 0, 0, 0,
  2.377197e-014, 1.803664e-014, 2.451693e-011, 3.347559e-011,
  0, 0, 0, 0,
  5.201021e-014, 1.850946e-014, 2.586179e-011, 4.587505e-011,
  0, 0, 0, 0,
  8.355272e-015, 3.019773e-014, 3.397689e-011, 5.05916e-011,
  0, 0, 0, 0,
  6.772167e-015, 1.335624e-014, 2.378947e-011, 3.573349e-011,
  0, 0, 0, 0,
  5.902117e-015, 1.542115e-014, 2.814413e-011, 5.010048e-011,
  0, 0, 0, 0,
  7.543607e-014, 1.404855e-014, 2.22021e-011, 3.196508e-011,
  0, 0, 0, 0,
  3.537094e-015, 7.551441e-015, 2.138361e-011, 3.655629e-011,
  0, 0, 0, 0,
  2.663662e-015, 2.658703e-015, 1.137079e-011, 1.297957e-011,
  0, 0, 0, 0,
  1.859426e-015, 4.369104e-015, 1.054473e-011, 1.373661e-011,
  0, 0, 0, 0,
  3.156845e-015, 4.787973e-015, 4.614613e-012, 8.293395e-012,
  0, 0, 0, 0,
  2.650043e-015, 4.628979e-015, 5.86769e-012, 9.206961e-012,
  0, 0, 0, 0,
  2.33386e-015, 4.988745e-015, 8.559323e-012, 1.138404e-011,
  0, 0, 0, 0,
  2.44409e-014, 1.186166e-014, 1.034253e-011, 1.646837e-011,
  0, 0, 0, 0,
  5.016386e-014, 9.027229e-015, 9.400958e-012, 1.574363e-011,
  0, 0, 0, 0,
  2.355766e-014, 1.21804e-014, 1.495627e-011, 1.988517e-011,
  0, 0, 0, 0,
  5.350324e-014, 2.425882e-014, 1.386488e-011, 3.217803e-011,
  0, 0, 0, 0,
  1.131611e-014, 9.090979e-015, 1.727666e-011, 3.325801e-011,
  0, 0, 0, 0,
  2.666703e-014, 7.014723e-015, 1.327705e-011, 2.503603e-011,
  0, 0, 0, 0,
  5.181454e-014, 1.076257e-014, 2.768647e-011, 3.995784e-011,
  0, 0, 0, 0,
  4.979759e-015, 1.012253e-014, 3.022972e-011, 5.243573e-011,
  0, 0, 0, 0,
  5.173585e-015, 5.274782e-015, 2.007099e-011, 3.865726e-011,
  0, 0, 0, 0,
  8.408627e-015, 6.538337e-015, 3.960193e-011, 6.838543e-011,
  0, 0, 0, 0,
  9.744602e-015, 1.902644e-014, 6.890152e-011, 9.882305e-011,
  0, 0, 0, 0,
  5.919176e-015, 4.157182e-015, 3.271483e-011, 5.001299e-011,
  0, 0, 0, 0,
  7.319242e-015, 4.515519e-015, 3.217646e-011, 5.303435e-011,
  0, 0, 0, 0,
  7.863234e-015, 1.356312e-014, 2.909359e-011, 4.763691e-011,
  0, 0, 0, 0,
  7.059571e-014, 1.665601e-014, 4.049052e-011, 6.902005e-011,
  0, 0, 0, 0,
  7.779022e-015, 1.34578e-014, 3.397416e-011, 4.847994e-011,
  0, 0, 0, 0,
  8.104565e-015, 2.04079e-014, 3.819334e-011, 5.234825e-011,
  0, 0, 0, 0,
  8.53538e-015, 2.714484e-014, 4.19579e-011, 7.158164e-011,
  0, 0, 0, 0,
  6.09478e-014, 2.780687e-014, 5.705254e-011, 7.872929e-011,
  0, 0, 0, 0,
  2.430419e-014, 3.669108e-014, 6.633966e-011, 9.819656e-011,
  0, 0, 0, 0,
  1.252115e-014, 2.778771e-014, 4.075152e-011, 6.457062e-011,
  0, 0, 0, 0,
  1.271018e-014, 4.011215e-014, 4.363424e-011, 8.419489e-011,
  0, 0, 0, 0,
  1.062293e-014, 3.557697e-014, 6.502257e-011, 1.070579e-010,
  0, 0, 0, 0,
  7.527572e-015, 2.159447e-014, 3.77937e-011, 6.298539e-011,
  0, 0, 0, 0,
  6.199682e-015, 2.00904e-014, 3.25495e-011, 5.581039e-011,
  0, 0, 0, 0,
  5.439801e-015, 1.495689e-014, 2.491731e-011, 4.467798e-011,
  0, 0, 0, 0,
  1.310949e-014, 1.574242e-014, 2.854567e-011, 4.724411e-011,
  0, 0, 0, 0,
  6.651799e-014, 1.190007e-014, 2.206067e-011, 3.644342e-011,
  0, 0, 0, 0,
  5.434992e-015, 6.069734e-015, 2.117525e-011, 3.433359e-011,
  0, 0, 0, 0,
  5.267136e-015, 6.572758e-015, 2.056752e-011, 3.719358e-011,
  0, 0, 0, 0,
  6.667092e-015, 1.374985e-014, 2.689279e-011, 4.692208e-011,
  0, 0, 0, 0,
  7.285765e-014, 1.311015e-014, 1.988754e-011, 3.27044e-011,
  0, 0, 0, 0,
  4.930548e-015, 1.053432e-014, 1.94865e-011, 3.563116e-011,
  0, 0, 0, 0,
  6.355671e-015, 1.538659e-014, 2.372223e-011, 4.717537e-011,
  0, 0, 0, 0,
  1.068305e-014, 3.261843e-014, 4.265099e-011, 7.51129e-011,
  0, 0, 0, 0,
  5.649437e-015, 1.784828e-014, 2.305965e-011, 4.19285e-011,
  0, 0, 0, 0,
  5.471759e-015, 1.288726e-014, 2.3547e-011, 4.222513e-011,
  0, 0, 0, 0,
  8.602876e-015, 3.777614e-014, 2.576277e-011, 5.45907e-011,
  0, 0, 0, 0,
  7.679823e-015, 3.461434e-014, 3.018136e-011, 4.363489e-011,
  0, 0, 0, 0,
  9.28672e-015, 2.474825e-014, 3.735936e-011, 5.561672e-011,
  0, 0, 0, 0,
  1.257057e-014, 2.928037e-014, 4.002735e-011, 7.288378e-011,
  0, 0, 0, 0,
  7.839629e-015, 1.788713e-014, 4.510618e-011, 7.457978e-011,
  0, 0, 0, 0,
  8.130725e-015, 1.815483e-014, 3.016831e-011, 4.893139e-011,
  0, 0, 0, 0,
  1.934505e-014, 2.235004e-014, 2.979059e-011, 4.537976e-011,
  0, 0, 0, 0,
  5.80943e-014, 3.383002e-014, 3.148363e-011, 5.276462e-011,
  0, 0, 0, 0,
  6.383289e-015, 2.218337e-014, 4.210747e-011, 6.62365e-011,
  0, 0, 0, 0,
  5.239644e-015, 1.910287e-014, 3.698836e-011, 5.945868e-011,
  0, 0, 0, 0,
  5.852183e-015, 1.756447e-014, 2.53583e-011, 4.071025e-011,
  0, 0, 0, 0,
  7.169293e-014, 1.706516e-014, 2.464903e-011, 5.012739e-011,
  0, 0, 0, 0,
  6.309398e-015, 1.564398e-014, 2.812715e-011, 4.845261e-011,
  0, 0, 0, 0,
  5.536074e-015, 3.023897e-014, 1.679257e-011, 3.89752e-011,
  0, 0, 0, 0,
  5.912807e-015, 2.207163e-014, 2.942337e-011, 4.687516e-011,
  0, 0, 0, 0,
  6.133327e-015, 2.431581e-014, 2.064464e-011, 4.097845e-011,
  0, 0, 0, 0,
  5.858645e-015, 2.105105e-014, 3.242772e-011, 5.558156e-011,
  0, 0, 0, 0,
  6.755029e-015, 2.467517e-014, 2.153209e-011, 4.041465e-011,
  0, 0, 0, 0,
  7.794296e-015, 2.576154e-014, 2.40724e-011, 4.845965e-011,
  0, 0, 0, 0,
  5.487244e-014, 2.856715e-014, 2.381537e-011, 4.295753e-011,
  0, 0, 0, 0,
  1.717567e-014, 2.375112e-014, 5.491096e-011, 9.03613e-011,
  0, 0, 0, 0,
  1.144141e-014, 2.369672e-014, 5.329196e-011, 7.988344e-011,
  0, 0, 0, 0,
  1.219703e-014, 2.775842e-014, 3.112727e-011, 4.929323e-011,
  0, 0, 0, 0,
  2.856988e-014, 2.145101e-014, 4.601537e-011, 7.361067e-011,
  0, 0, 0, 0,
  5.212009e-014, 2.407267e-014, 4.649561e-011, 8.606166e-011,
  0, 0, 0, 0,
  6.993725e-015, 2.230979e-014, 4.850972e-011, 7.501971e-011,
  0, 0, 0, 0,
  9.305719e-015, 2.340233e-014, 3.428885e-011, 6.11527e-011,
  0, 0, 0, 0,
  6.95679e-015, 2.511334e-014, 3.482381e-011, 6.097226e-011,
  0, 0, 0, 0,
  1.078247e-014, 1.531917e-014, 3.764931e-011, 5.243316e-011,
  0, 0, 0, 0,
  5.816331e-015, 1.228085e-014, 2.220717e-011, 3.861173e-011,
  0, 0, 0, 0,
  6.719348e-015, 2.177303e-014, 3.20521e-011, 6.023666e-011,
  0, 0, 0, 0,
  9.020083e-015, 1.732972e-014, 6.455059e-011, 9.917659e-011,
  0, 0, 0, 0,
  7.041342e-014, 2.276157e-014, 2.769778e-011, 4.454117e-011,
  0, 0, 0, 0,
  5.011861e-015, 2.199856e-014, 2.806703e-011, 5.718898e-011,
  0, 0, 0, 0,
  5.209815e-015, 1.662846e-014, 2.775545e-011, 3.960311e-011,
  0, 0, 0, 0,
  6.93005e-015, 1.924466e-014, 3.575332e-011, 5.863999e-011,
  0, 0, 0, 0,
  6.71141e-014, 2.322528e-014, 4.028305e-011, 5.312392e-011,
  0, 0, 0, 0,
  1.385109e-014, 1.854359e-014, 2.400239e-011, 4.696542e-011,
  0, 0, 0, 0,
  5.922172e-015, 1.575324e-014, 2.306053e-011, 3.79819e-011,
  0, 0, 0, 0,
  6.894043e-015, 1.604298e-014, 3.434297e-011, 5.353013e-011,
  0, 0, 0, 0,
  8.64299e-015, 2.526003e-014, 4.275601e-011, 7.127171e-011,
  0, 0, 0, 0,
  8.637282e-015, 2.8609e-014, 2.963539e-011, 4.340763e-011,
  0, 0, 0, 0,
  6.999613e-015, 1.313306e-014, 3.434819e-011, 5.523211e-011,
  0, 0, 0, 0,
  1.266247e-014, 1.71776e-014, 3.882252e-011, 6.92767e-011,
  0, 0, 0, 0,
  1.224711e-014, 2.322797e-014, 3.841845e-011, 6.834043e-011,
  0, 0, 0, 0,
  2.829849e-014, 1.994156e-014, 3.964352e-011, 6.038567e-011,
  0, 0, 0, 0,
  1.627715e-014, 5.757188e-014, 4.920308e-011, 9.678244e-011,
  0, 0, 0, 0,
  1.028776e-014, 3.638157e-014, 4.177197e-011, 7.087256e-011,
  0, 0, 0, 0,
  1.334887e-014, 2.537298e-014, 5.418754e-011, 1.029249e-010,
  0, 0, 0, 0,
  2.296315e-015, 2.140239e-015, 4.713614e-012, 4.30258e-012,
  0, 0, 0, 0,
  1.805057e-014, 3.942538e-015, 3.379548e-011, 2.804788e-011,
  0, 0, 0, 0,
  6.018853e-014, 9.574611e-015, 4.473305e-012, 4.118757e-012,
  0, 0, 0, 0,
  8.331629e-015, 5.493666e-015, 1.15688e-011, 1.827069e-011,
  0, 0, 0, 0,
  4.061615e-015, 3.460445e-015, 3.858132e-012, 4.644609e-012,
  0, 0, 0, 0,
  2.980208e-015, 3.562851e-015, 1.407646e-011, 1.765816e-011,
  0, 0, 0, 0,
  7.676737e-014, 1.233966e-014, 6.440058e-012, 6.924649e-012,
  0, 0, 0, 0,
  2.124298e-015, 3.443239e-015, 6.018621e-012, 8.382003e-012,
  0, 0, 0, 0,
  1.489603e-014, 3.287195e-015, 9.217513e-012, 7.584859e-012,
  0, 0, 0, 0,
  1.719269e-014, 8.1893e-014, 7.306405e-012, 5.975675e-012,
  0, 0, 0, 0,
  7.464245e-014, 1.565288e-014, 3.709855e-012, 4.98968e-012,
  0, 0, 0, 0,
  8.723331e-015, 2.181554e-015, 3.125511e-012, 3.41262e-012,
  0, 0, 0, 0,
  2.603497e-015, 1.707906e-015, 4.580465e-012, 5.805909e-012,
  0, 0, 0, 0,
  2.810669e-015, 2.140436e-015, 5.902263e-012, 7.003945e-012,
  0, 0, 0, 0,
  3.339239e-015, 2.252277e-015, 3.487683e-012, 5.605437e-012,
  0, 0, 0, 0,
  2.884083e-015, 2.131174e-015, 6.189032e-012, 7.515436e-012,
  0, 0, 0, 0,
  5.526289e-015, 2.382516e-015, 1.01135e-011, 1.598296e-011,
  0, 0, 0, 0,
  2.146031e-015, 2.565317e-015, 3.756274e-012, 5.099416e-012,
  0, 0, 0, 0,
  3.08268e-015, 6.296484e-015, 3.871342e-012, 4.709833e-012,
  0, 0, 0, 0,
  3.385564e-015, 2.929559e-015, 4.352071e-012, 4.185214e-012,
  0, 0, 0, 0,
  2.537798e-015, 3.047658e-015, 6.656042e-012, 7.875501e-012,
  0, 0, 0, 0,
  2.659522e-015, 1.900168e-015, 5.662657e-012, 5.637871e-012,
  0, 0, 0, 0,
  8.329248e-015, 2.162366e-015, 5.74961e-012, 8.362803e-012,
  0, 0, 0, 0,
  6.919775e-014, 1.12215e-014, 4.556714e-012, 6.454828e-012,
  0, 0, 0, 0,
  3.446595e-015, 1.606567e-014, 6.211386e-012, 9.565985e-012,
  0, 0, 0, 0,
  1.99654e-015, 8.102697e-015, 5.067453e-012, 6.432759e-012,
  0, 0, 0, 0,
  3.923018e-015, 7.978844e-015, 4.622267e-012, 8.126642e-012,
  0, 0, 0, 0,
  8.364249e-014, 1.318416e-014, 1.390002e-011, 1.813914e-011,
  0, 0, 0, 0,
  3.51983e-015, 2.643899e-015, 7.647187e-012, 1.077582e-011,
  0, 0, 0, 0,
  3.117762e-015, 3.817814e-015, 5.958885e-012, 7.443281e-012,
  0, 0, 0, 0,
  2.190614e-015, 2.045965e-015, 2.516401e-012, 3.312606e-012,
  0, 0, 0, 0,
  4.566801e-015, 1.62991e-015, 1.417446e-011, 6.678205e-011,
  0, 0, 0, 0,
  2.995108e-015, 1.912099e-015, 4.084243e-012, 4.350345e-012,
  0, 0, 0, 0,
  1.164823e-014, 2.50308e-015, 4.053583e-012, 5.937005e-012,
  0, 0, 0, 0,
  3.530969e-015, 3.365704e-015, 4.845906e-012, 5.154469e-012,
  0, 0, 0, 0,
  3.99611e-014, 7.622588e-015, 5.94212e-012, 8.028905e-012,
  0, 0, 0, 0,
  4.801534e-014, 7.710021e-015, 5.566144e-012, 6.159776e-012,
  0, 0, 0, 0,
  2.315102e-015, 1.708889e-015, 3.624354e-012, 5.120573e-012,
  0, 0, 0, 0,
  6.718464e-015, 2.378307e-015, 3.093115e-012, 3.054866e-012,
  0, 0, 0, 0,
  1.280113e-014, 2.641712e-015, 2.548623e-012, 3.264391e-012,
  0, 0, 0, 0,
  7.479523e-014, 1.178305e-014, 2.593598e-012, 4.141742e-012,
  0, 0, 0, 0,
  6.25342e-015, 2.213181e-015, 5.706918e-012, 7.278376e-012,
  0, 0, 0, 0,
  2.883796e-015, 2.7376e-015, 3.657321e-012, 5.549194e-012,
  0, 0, 0, 0,
  2.389585e-015, 2.194245e-015, 4.821426e-012, 4.041733e-012,
  0, 0, 0, 0,
  8.243628e-014, 1.274825e-014, 3.676177e-012, 4.023856e-012,
  0, 0, 0, 0,
  2.9366e-015, 2.156887e-015, 3.841307e-012, 5.39413e-012,
  0, 0, 0, 0,
  2.759279e-015, 3.419707e-015, 4.908453e-012, 1.099993e-011,
  0, 0, 0, 0,
  1.839294e-015, 5.655851e-015, 3.370641e-012, 4.302192e-012,
  0, 0, 0, 0,
  7.395531e-014, 2.789658e-014, 4.362919e-012, 6.485754e-012,
  0, 0, 0, 0,
  1.015208e-014, 3.329914e-015, 1.771197e-011, 1.853035e-011,
  0, 0, 0, 0,
  2.576944e-015, 4.24471e-015, 2.58058e-012, 3.268354e-012,
  0, 0, 0, 0,
  2.359716e-015, 4.490712e-015, 3.205151e-012, 3.393012e-012,
  0, 0, 0, 0,
  4.232185e-014, 7.089374e-015, 3.50939e-012, 4.346806e-012,
  0, 0, 0, 0,
  3.228731e-014, 7.721449e-015, 4.614612e-012, 5.245509e-012,
  0, 0, 0, 0,
  1.659213e-015, 1.62022e-015, 4.126918e-012, 3.21805e-012,
  0, 0, 0, 0,
  2.853616e-015, 1.856811e-015, 2.944687e-012, 3.380744e-012,
  0, 0, 0, 0,
  2.289328e-014, 4.301831e-015, 4.159981e-012, 4.23107e-012,
  0, 0, 0, 0,
  5.806216e-014, 9.26752e-015, 5.205937e-012, 4.817703e-012,
  0, 0, 0, 0,
  2.350469e-015, 2.724283e-015, 3.71864e-012, 3.795331e-012,
  0, 0, 0, 0,
  1.431786e-015, 1.951479e-015, 2.816015e-012, 2.835821e-012,
  0, 0, 0, 0,
  2.388933e-015, 2.637325e-015, 2.94145e-012, 3.059159e-012,
  0, 0, 0, 0,
  2.454839e-015, 2.496439e-015, 2.813962e-012, 3.007228e-012,
  0, 0, 0, 0,
  2.519888e-015, 1.372271e-015, 2.453565e-012, 2.813742e-012,
  0, 0, 0, 0,
  1.665693e-015, 2.064233e-015, 2.257291e-012, 2.697445e-012,
  0, 0, 0, 0,
  2.489905e-015, 3.289734e-015, 2.806501e-012, 2.334851e-012,
  0, 0, 0, 0,
  7.512796e-014, 1.231897e-014, 4.878147e-012, 6.285728e-012,
  0, 0, 0, 0,
  3.555422e-015, 2.134835e-015, 3.490133e-012, 3.652648e-012,
  0, 0, 0, 0,
  2.078852e-015, 5.447156e-015, 5.572764e-012, 9.460343e-012,
  0, 0, 0, 0,
  3.34064e-015, 5.771174e-015, 7.16087e-012, 1.204253e-011,
  0, 0, 0, 0,
  5.87359e-014, 9.599612e-015, 3.435178e-012, 3.752625e-012,
  0, 0, 0, 0,
  1.751282e-014, 3.391474e-015, 4.40837e-012, 4.96968e-012,
  0, 0, 0, 0,
  3.166902e-015, 2.960001e-015, 1.324103e-011, 1.478652e-011,
  0, 0, 0, 0,
  2.452969e-015, 2.527142e-015, 3.187493e-012, 4.701015e-012,
  0, 0, 0, 0,
  3.324302e-014, 5.62355e-015, 2.53242e-012, 3.495847e-012,
  0, 0, 0, 0,
  4.893642e-014, 7.655484e-015, 2.141164e-012, 2.546707e-012,
  0, 0, 0, 0,
  2.426244e-015, 2.886317e-015, 3.332044e-012, 4.150987e-012,
  0, 0, 0, 0,
  4.256986e-015, 1.986079e-015, 3.823738e-012, 4.829457e-012,
  0, 0, 0, 0,
  4.420455e-015, 2.554161e-015, 3.915239e-012, 5.251384e-012,
  0, 0, 0, 0,
  5.07265e-015, 4.003098e-015, 4.779155e-012, 6.630454e-012,
  0, 0, 0, 0,
  3.48957e-015, 4.187397e-015, 4.850031e-012, 8.676458e-012,
  0, 0, 0, 0,
  3.358113e-015, 3.286174e-015, 7.544434e-012, 7.096613e-012,
  0, 0, 0, 0,
  3.856433e-015, 4.593399e-015, 9.855886e-012, 1.404415e-011,
  0, 0, 0, 0,
  8.284991e-014, 1.343466e-014, 5.690364e-012, 7.268935e-012,
  0, 0, 0, 0,
  2.925381e-015, 4.139134e-015, 1.511967e-011, 2.224288e-011,
  0, 0, 0, 0,
  3.650447e-015, 5.893077e-015, 6.596062e-012, 1.204205e-011,
  0, 0, 0, 0,
  3.454949e-015, 5.296788e-015, 1.313038e-011, 1.619511e-011,
  0, 0, 0, 0,
  6.933463e-014, 1.149339e-014, 5.047483e-012, 5.741168e-012,
  0, 0, 0, 0,
  1.024697e-014, 4.248284e-015, 5.688667e-012, 8.482828e-012,
  0, 0, 0, 0,
  4.05543e-015, 4.166807e-015, 7.015241e-012, 1.00529e-011,
  0, 0, 0, 0,
  3.97156e-015, 1.339725e-014, 1.324772e-011, 1.743988e-011,
  0, 0, 0, 0,
  5.170169e-014, 1.138475e-014, 6.308087e-012, 1.171897e-011,
  0, 0, 0, 0,
  3.195322e-014, 7.29786e-015, 9.916158e-012, 1.706876e-011,
  0, 0, 0, 0,
  4.224087e-015, 5.386858e-015, 9.108954e-012, 1.312456e-011,
  0, 0, 0, 0,
  5.61352e-015, 3.673866e-015, 1.510293e-011, 1.78422e-011,
  0, 0, 0, 0,
  7.857117e-015, 4.151829e-015, 6.118117e-012, 9.860689e-012,
  0, 0, 0, 0,
  2.227641e-015, 3.926499e-015, 6.385127e-012, 7.501028e-012,
  0, 0, 0, 0,
  2.750478e-015, 3.695494e-015, 5.210794e-012, 6.259508e-012,
  0, 0, 0, 0,
  2.949806e-015, 3.111887e-015, 4.93119e-012, 4.874772e-012,
  0, 0, 0, 0,
  3.75123e-015, 3.588011e-015, 4.498005e-012, 8.492012e-012,
  0, 0, 0, 0,
  2.026827e-015, 3.168337e-015, 4.310664e-012, 4.197401e-012,
  0, 0, 0, 0,
  1.66558e-015, 1.879708e-015, 3.621318e-012, 3.542712e-012,
  0, 0, 0, 0,
  2.889425e-015, 3.768857e-015, 3.227801e-012, 3.23623e-012,
  0, 0, 0, 0,
  6.424371e-014, 1.006175e-014, 1.246099e-011, 1.516753e-011,
  0, 0, 0, 0,
  1.01517e-014, 3.552271e-015, 3.431188e-011, 4.091599e-011,
  0, 0, 0, 0,
  9.654814e-015, 5.777749e-015, 2.768526e-011, 4.205908e-011,
  0, 0, 0, 0,
  6.162957e-014, 1.485304e-014, 6.450185e-011, 1.015299e-010,
  0, 0, 0, 0,
  6.226681e-015, 4.701328e-015, 6.631239e-012, 8.037447e-012,
  0, 0, 0, 0,
  9.616407e-015, 4.906598e-015, 5.020157e-012, 4.460788e-012,
  0, 0, 0, 0,
  1.103604e-014, 6.173925e-015, 2.198729e-011, 3.412027e-011,
  0, 0, 0, 0,
  2.2188e-014, 6.577447e-015, 4.794688e-012, 1.031524e-011,
  0, 0, 0, 0,
  2.343441e-014, 8.69168e-015, 5.306822e-012, 7.683492e-012,
  0, 0, 0, 0,
  2.533005e-014, 6.710001e-015, 3.434924e-012, 5.840223e-012,
  0, 0, 0, 0,
  4.195387e-014, 1.210819e-014, 5.41034e-012, 7.113533e-012,
  0, 0, 0, 0,
  6.318256e-014, 1.408184e-014, 4.465248e-012, 1.315109e-011,
  0, 0, 0, 0,
  9.354853e-014, 1.942888e-014, 7.829361e-012, 1.770826e-011,
  0, 0, 0, 0,
  5.583113e-014, 1.337782e-014, 1.712187e-011, 2.056277e-011,
  0, 0, 0, 0,
  9.005372e-014, 1.861246e-014, 4.782415e-012, 1.360764e-011,
  0, 0, 0, 0,
  1.09229e-013, 3.334349e-014, 5.154353e-012, 1.586073e-011,
  0, 0, 0, 0,
  1.469347e-013, 4.391347e-014, 5.816703e-012, 1.896999e-011,
  0, 0, 0, 0,
  3.705526e-013, 6.834171e-014, 1.261925e-011, 6.230972e-011,
  0, 0, 0, 0,
  3.140409e-013, 7.565096e-014, 8.953473e-012, 3.730974e-011,
  0, 0, 0, 0,
  7.075085e-013, 1.350797e-013, 2.22672e-011, 9.747807e-011,
  0, 0, 0, 0,
  7.87735e-013, 1.657411e-013, 2.358667e-011, 1.043134e-010,
  0, 0, 0, 0,
  1.263043e-012, 2.787747e-013, 4.11498e-011, 1.805874e-010,
  0, 0, 0, 0,
  1.639463e-012, 3.481729e-013, 1.001397e-010, 4.143854e-010,
  0, 0, 0, 0,
  2.522678e-012, 6.100835e-013, 9.231016e-011, 4.010378e-010,
  0, 0, 0, 0,
  3.789811e-012, 1.089867e-012, 1.815436e-010, 6.885553e-010,
  0, 0, 0, 0,
  6.229049e-012, 2.152581e-012, 6.609842e-010, 1.708895e-009,
  0, 0, 0, 0,
  1.346614e-011, 4.26248e-012, 1.378668e-009, 7.013998e-009,
  0, 0, 0, 0,
  1.550391e-011, 4.415109e-012, 9.895541e-010, 3.428355e-009,
  0, 0, 0, 0,
  8.347125e-012, 3.199094e-012, 8.81803e-010, 2.559096e-009,
  0, 0, 0, 0,
  1.275366e-011, 3.411751e-012, 8.8211e-010, 2.697972e-009,
  0, 0, 0, 0,
  1.345067e-011, 4.625157e-012, 9.17812e-010, 3.549933e-009,
  0, 0, 0, 0,
  4.05514e-012, 2.170539e-012, 3.619948e-010, 1.381968e-009,
  0, 0, 0, 0,
  3.434263e-012, 7.187248e-013, 1.324232e-010, 5.794327e-010,
  0, 0, 0, 0,
  1.89742e-012, 5.721626e-013, 6.90968e-011, 2.979041e-010,
  0, 0, 0, 0,
  1.543477e-012, 3.67044e-013, 5.64463e-011, 2.272924e-010,
  0, 0, 0, 0,
  1.080035e-012, 3.621159e-013, 4.311359e-011, 1.345528e-010,
  0, 0, 0, 0,
  4.958581e-013, 2.307136e-013, 3.457533e-011, 1.286836e-010,
  0, 0, 0, 0,
  3.333436e-013, 2.266585e-013, 1.869643e-011, 5.693967e-011,
  0, 0, 0, 0,
  2.762448e-013, 1.736354e-013, 2.050846e-011, 5.284094e-011,
  0, 0, 0, 0,
  1.974167e-013, 1.245317e-013, 2.24982e-011, 8.008409e-011,
  0, 0, 0, 0,
  1.618312e-013, 3.885243e-014, 1.191992e-011, 2.063278e-011,
  0, 0, 0, 0,
  9.591393e-014, 2.654889e-014, 1.323278e-011, 3.02422e-011,
  0, 0, 0, 0,
  1.443092e-013, 3.707249e-014, 8.56023e-012, 2.536732e-011,
  0, 0, 0, 0,
  7.547712e-014, 1.127176e-013, 1.853988e-011, 6.345918e-011,
  0, 0, 0, 0,
  4.240207e-014, 1.793929e-014, 5.459121e-012, 9.480214e-012,
  0, 0, 0, 0,
  2.997196e-014, 1.28337e-014, 7.547034e-012, 1.131869e-011,
  0, 0, 0, 0,
  2.477684e-014, 2.64202e-014, 1.47533e-011, 3.179043e-011,
  0, 0, 0, 0,
  3.31725e-014, 2.280613e-014, 9.765303e-012, 2.472102e-011,
  0, 0, 0, 0,
  3.278889e-014, 4.658546e-014, 3.603829e-011, 6.714496e-011,
  0, 0, 0, 0,
  2.473e-014, 5.929109e-014, 3.467776e-011, 7.43564e-011,
  0, 0, 0, 0,
  3.989574e-014, 2.358646e-013, 4.278282e-011, 1.525727e-010,
  0, 0, 0, 0,
  7.480693e-014, 6.32335e-014, 2.95741e-011, 7.250266e-011,
  0, 0, 0, 0,
  1.77959e-014, 7.471098e-014, 2.515579e-011, 5.665419e-011,
  0, 0, 0, 0,
  1.169029e-014, 4.134316e-014, 1.514575e-011, 2.996072e-011,
  0, 0, 0, 0,
  5.664516e-015, 2.145863e-014, 1.35475e-011, 2.196571e-011,
  0, 0, 0, 0,
  8.453062e-015, 4.541094e-014, 2.137374e-011, 3.555362e-011,
  0, 0, 0, 0,
  3.869206e-015, 1.215128e-014, 1.778139e-011, 3.329529e-011,
  0, 0, 0, 0,
  4.511745e-015, 7.312758e-015, 1.875721e-011, 2.061495e-011,
  0, 0, 0, 0,
  4.756241e-015, 9.167189e-015, 6.228115e-012, 8.149386e-012,
  0, 0, 0, 0,
  7.511404e-015, 4.653599e-014, 1.637352e-011, 3.712355e-011,
  0, 0, 0, 0,
  4.351295e-015, 1.022333e-014, 4.864483e-012, 8.876145e-012,
  0, 0, 0, 0,
  4.88858e-015, 1.241085e-014, 6.383334e-012, 1.034267e-011,
  0, 0, 0, 0,
  3.896386e-015, 1.942437e-014, 7.473815e-012, 1.717816e-011,
  0, 0, 0, 0,
  1.469122e-014, 1.524222e-014, 1.012877e-011, 2.35476e-011,
  0, 0, 0, 0,
  4.031739e-015, 1.829719e-014, 8.446717e-012, 1.501744e-011,
  0, 0, 0, 0,
  9.557395e-015, 5.072195e-014, 2.876432e-011, 7.010702e-011,
  0, 0, 0, 0,
  1.498195e-014, 7.911788e-014, 2.153066e-011, 5.478848e-011,
  0, 0, 0, 0,
  4.340349e-014, 2.710837e-013, 4.328359e-011, 1.447829e-010,
  0, 0, 0, 0,
  7.920119e-014, 7.373458e-014, 3.701986e-011, 7.188244e-011,
  0, 0, 0, 0,
  2.438347e-014, 1.511913e-013, 7.269262e-011, 1.639392e-010,
  0, 0, 0, 0,
  2.371784e-014, 1.485505e-013, 4.810606e-011, 1.138441e-010,
  0, 0, 0, 0,
  9.608328e-015, 5.025582e-014, 2.012895e-011, 4.146974e-011,
  0, 0, 0, 0,
  6.452186e-014, 7.395863e-014, 2.549657e-011, 7.260122e-011,
  0, 0, 0, 0,
  1.192551e-014, 4.108653e-014, 3.035406e-011, 6.465061e-011,
  0, 0, 0, 0,
  3.634975e-015, 1.355913e-014, 7.139081e-012, 1.342119e-011,
  0, 0, 0, 0,
  1.535478e-014, 9.711362e-014, 2.096925e-011, 5.76916e-011,
  0, 0, 0, 0,
  4.914839e-014, 9.624609e-014, 1.538363e-011, 5.428239e-011,
  0, 0, 0, 0,
  2.959242e-014, 2.383185e-014, 1.006008e-011, 1.808972e-011,
  0, 0, 0, 0,
  1.694969e-014, 9.804427e-014, 2.212143e-011, 6.461246e-011,
  0, 0, 0, 0,
  1.010341e-014, 4.700868e-014, 1.940405e-011, 4.548447e-011,
  0, 0, 0, 0,
  2.589367e-014, 1.609299e-013, 3.723727e-011, 1.140031e-010,
  0, 0, 0, 0,
  1.202593e-014, 6.027053e-014, 1.966617e-011, 4.832375e-011,
  0, 0, 0, 0,
  3.683279e-014, 2.345588e-013, 3.927726e-011, 1.25163e-010,
  0, 0, 0, 0,
  2.161013e-014, 1.343004e-013, 4.464999e-011, 1.147202e-010,
  0, 0, 0, 0,
  3.742635e-014, 2.402497e-013, 7.559631e-011, 1.953644e-010,
  0, 0, 0, 0,
  7.697508e-014, 6.592413e-014, 4.019162e-011, 8.293208e-011,
  0, 0, 0, 0,
  2.171244e-014, 1.357059e-013, 4.481401e-011, 1.1758e-010,
  0, 0, 0, 0,
  2.084501e-014, 1.24876e-013, 3.864575e-011, 9.974487e-011,
  0, 0, 0, 0,
  3.170293e-014, 2.019383e-013, 4.810019e-011, 1.469543e-010,
  0, 0, 0, 0,
  6.974964e-014, 7.69915e-014, 1.769147e-011, 5.473739e-011,
  0, 0, 0, 0,
  5.831959e-015, 2.389421e-014, 2.079774e-011, 4.067715e-011,
  0, 0, 0, 0,
  6.224341e-015, 2.094517e-014, 1.475938e-011, 2.412055e-011,
  0, 0, 0, 0,
  8.739232e-015, 5.362328e-014, 1.01327e-011, 3.347323e-011,
  0, 0, 0, 0,
  5.814548e-014, 2.000596e-014, 7.75635e-012, 1.355508e-011,
  0, 0, 0, 0,
  2.042358e-014, 7.091512e-015, 5.404996e-012, 7.140464e-012,
  0, 0, 0, 0,
  4.149794e-015, 1.411141e-014, 1.131254e-011, 1.744282e-011,
  0, 0, 0, 0,
  3.721893e-015, 1.624883e-014, 5.825556e-012, 1.329873e-011,
  0, 0, 0, 0,
  5.049325e-015, 2.010902e-014, 1.676974e-011, 3.864832e-011,
  0, 0, 0, 0,
  4.155029e-015, 2.430926e-014, 1.454702e-011, 2.995756e-011,
  0, 0, 0, 0,
  5.345436e-015, 2.430894e-014, 1.460415e-011, 3.029495e-011,
  0, 0, 0, 0,
  4.085006e-015, 1.755822e-014, 1.482987e-011, 3.292213e-011,
  0, 0, 0, 0,
  2.094579e-014, 1.035024e-013, 1.948369e-011, 6.092279e-011,
  0, 0, 0, 0,
  7.979816e-014, 1.391871e-013, 2.51426e-011, 8.713531e-011,
  0, 0, 0, 0,
  1.321608e-014, 7.821275e-014, 3.466312e-011, 7.797545e-011,
  0, 0, 0, 0,
  4.462503e-014, 2.866955e-013, 8.150113e-011, 2.138137e-010,
  0, 0, 0, 0,
  3.619115e-014, 2.189727e-013, 5.16162e-011, 1.270434e-010,
  0, 0, 0, 0,
  8.447113e-014, 2.574785e-013, 7.678932e-011, 2.046317e-010,
  0, 0, 0, 0,
  2.628135e-014, 1.63228e-013, 7.791942e-011, 1.684114e-010,
  0, 0, 0, 0,
  6.718976e-014, 4.269994e-013, 1.322886e-010, 3.366874e-010,
  0, 0, 0, 0,
  3.012561e-014, 1.79629e-013, 7.015256e-011, 1.505844e-010,
  0, 0, 0, 0,
  7.711221e-014, 1.213629e-013, 8.846384e-011, 1.633096e-010,
  0, 0, 0, 0,
  2.768997e-014, 1.010794e-013, 5.064403e-011, 9.054641e-011,
  0, 0, 0, 0,
  1.928088e-014, 1.072623e-013, 8.826138e-011, 1.511651e-010,
  0, 0, 0, 0,
  2.396442e-014, 8.350104e-014, 6.777197e-011, 1.165562e-010,
  0, 0, 0, 0,
  5.80248e-014, 1.958149e-013, 1.803343e-010, 2.605496e-010,
  0, 0, 0, 0,
  3.808345e-014, 1.129402e-013, 7.736076e-011, 1.013934e-010,
  0, 0, 0, 0,
  4.009265e-014, 1.752329e-013, 9.146425e-011, 1.632509e-010,
  0, 0, 0, 0,
  3.834661e-014, 2.344275e-013, 8.52446e-011, 1.992105e-010,
  0, 0, 0, 0,
  2.655871e-014, 8.069686e-014, 5.258092e-011, 8.463974e-011,
  0, 0, 0, 0,
  5.661078e-014, 8.889177e-014, 6.049802e-011, 1.157049e-010,
  0, 0, 0, 0,
  2.698515e-014, 1.444619e-013, 7.139022e-011, 1.335436e-010,
  0, 0, 0, 0,
  1.482281e-014, 2.726759e-014, 3.592792e-011, 5.821132e-011,
  0, 0, 0, 0,
  8.147887e-015, 1.804222e-014, 1.883239e-011, 2.862608e-011,
  0, 0, 0, 0,
  7.059085e-014, 1.770355e-014, 3.044663e-011, 4.209669e-011,
  0, 0, 0, 0,
  8.224287e-015, 1.039498e-014, 1.718789e-011, 2.731046e-011,
  0, 0, 0, 0,
  6.405687e-015, 3.318725e-015, 8.888347e-012, 1.512485e-011,
  0, 0, 0, 0,
  2.862379e-015, 4.253142e-015, 9.824354e-012, 1.522803e-011,
  0, 0, 0, 0,
  3.84956e-015, 3.471863e-015, 7.031956e-012, 9.783222e-012,
  0, 0, 0, 0,
  3.76881e-015, 7.355156e-015, 8.527716e-012, 1.261293e-011,
  0, 0, 0, 0,
  3.982341e-015, 5.160779e-015, 4.615998e-012, 6.47451e-012,
  0, 0, 0, 0,
  1.720648e-014, 1.048705e-014, 4.985427e-012, 6.750049e-012,
  0, 0, 0, 0,
  5.097822e-014, 1.387291e-014, 1.024133e-011, 2.033293e-011,
  0, 0, 0, 0,
  2.478269e-014, 2.806249e-014, 2.166203e-011, 4.203344e-011,
  0, 0, 0, 0,
  4.947526e-014, 9.700216e-014, 4.472165e-011, 8.769756e-011,
  0, 0, 0, 0,
  1.002723e-014, 8.857817e-015, 1.905292e-011, 3.180408e-011,
  0, 0, 0, 0,
  2.764318e-014, 8.164543e-015, 9.383471e-012, 1.793494e-011,
  0, 0, 0, 0,
  5.317648e-014, 1.516824e-014, 1.974245e-011, 2.823548e-011,
  0, 0, 0, 0,
  1.024216e-014, 2.138034e-014, 3.511125e-011, 3.675847e-011,
  0, 0, 0, 0,
  9.02848e-015, 7.807801e-015, 5.241861e-011, 8.794992e-011,
  0, 0, 0, 0,
  1.540699e-014, 1.658617e-014, 4.794629e-011, 7.095178e-011,
  0, 0, 0, 0,
  2.043709e-014, 5.065922e-014, 2.113142e-010, 2.818193e-010,
  0, 0, 0, 0,
  1.638315e-014, 1.199306e-014, 5.605968e-011, 7.65474e-011,
  0, 0, 0, 0,
  1.463032e-014, 1.055817e-014, 5.763777e-011, 9.436258e-011,
  0, 0, 0, 0,
  2.399705e-014, 1.259873e-014, 1.002238e-010, 1.466241e-010,
  0, 0, 0, 0,
  7.940739e-014, 2.251661e-014, 8.004021e-011, 1.341699e-010,
  0, 0, 0, 0,
  1.790201e-014, 2.688273e-014, 7.090765e-011, 1.289663e-010,
  0, 0, 0, 0,
  2.469068e-014, 4.746851e-014, 6.626703e-011, 1.107465e-010,
  0, 0, 0, 0,
  2.166642e-014, 1.051115e-013, 4.586133e-011, 7.546512e-011,
  0, 0, 0, 0,
  6.956257e-014, 1.262048e-013, 1.010626e-010, 1.5723e-010,
  0, 0, 0, 0,
  3.252428e-014, 1.363283e-013, 8.979185e-011, 1.525585e-010,
  0, 0, 0, 0,
  2.991415e-014, 1.202103e-013, 1.243303e-010, 1.93338e-010,
  0, 0, 0, 0,
  2.956952e-014, 1.647491e-013, 1.170254e-010, 1.828016e-010,
  0, 0, 0, 0,
  2.248217e-014, 4.987854e-014, 2.038473e-010, 2.860766e-010,
  0, 0, 0, 0,
  2.36084e-014, 7.210365e-014, 6.920065e-011, 1.14996e-010,
  0, 0, 0, 0,
  2.587104e-014, 1.071426e-013, 6.34397e-011, 1.400259e-010,
  0, 0, 0, 0,
  1.191736e-014, 2.480658e-014, 2.486015e-011, 3.529862e-011,
  0, 0, 0, 0,
  1.677313e-014, 1.973643e-014, 4.500062e-011, 6.626272e-011,
  0, 0, 0, 0,
  6.445372e-014, 1.468188e-014, 2.726e-011, 4.50515e-011,
  0, 0, 0, 0,
  8.653143e-015, 1.237359e-014, 2.578919e-011, 4.143127e-011,
  0, 0, 0, 0,
  7.539696e-015, 1.370311e-014, 2.134038e-011, 3.523161e-011,
  0, 0, 0, 0,
  9.720074e-015, 1.176057e-014, 2.846806e-011, 3.889291e-011,
  0, 0, 0, 0,
  7.382411e-014, 1.570848e-014, 2.208382e-011, 3.9226e-011,
  0, 0, 0, 0,
  5.784036e-015, 1.21831e-014, 1.383268e-011, 2.126659e-011,
  0, 0, 0, 0,
  1.370234e-014, 6.760935e-014, 5.04924e-011, 7.364283e-011,
  0, 0, 0, 0,
  4.928151e-014, 2.924714e-013, 1.19507e-010, 2.514296e-010,
  0, 0, 0, 0,
  1.882803e-014, 4.180626e-014, 3.970646e-011, 7.828185e-011,
  0, 0, 0, 0,
  1.269561e-014, 5.25047e-014, 4.384685e-011, 6.74365e-011,
  0, 0, 0, 0,
  2.763639e-014, 1.700917e-013, 4.118244e-011, 9.935715e-011,
  0, 0, 0, 0,
  3.236143e-014, 1.955467e-013, 6.972669e-011, 1.578091e-010,
  0, 0, 0, 0,
  2.826334e-014, 1.374159e-013, 5.800075e-011, 1.358337e-010,
  0, 0, 0, 0,
  2.57172e-014, 1.298714e-013, 4.564802e-011, 9.723108e-011,
  0, 0, 0, 0,
  2.403527e-014, 8.446392e-014, 7.536487e-011, 1.213791e-010,
  0, 0, 0, 0,
  1.659158e-014, 3.581074e-014, 4.034097e-011, 7.531611e-011,
  0, 0, 0, 0,
  2.180756e-014, 6.541028e-014, 5.704979e-011, 9.740959e-011,
  0, 0, 0, 0,
  6.062302e-014, 1.319827e-013, 6.707836e-011, 1.181778e-010,
  0, 0, 0, 0,
  1.856399e-014, 7.483661e-014, 4.726741e-011, 9.330335e-011,
  0, 0, 0, 0,
  1.58059e-014, 3.945363e-014, 5.291633e-011, 8.94582e-011,
  0, 0, 0, 0,
  2.162288e-014, 9.233503e-014, 4.510972e-011, 9.309565e-011,
  0, 0, 0, 0,
  7.867507e-014, 2.652716e-014, 2.720651e-011, 4.343275e-011,
  0, 0, 0, 0,
  1.446102e-014, 2.907802e-014, 4.121118e-011, 6.851786e-011,
  0, 0, 0, 0,
  2.596022e-014, 1.617775e-013, 2.930763e-011, 8.967303e-011,
  0, 0, 0, 0,
  2.676643e-014, 1.632023e-013, 4.799228e-011, 1.311501e-010,
  0, 0, 0, 0,
  1.614481e-014, 7.824432e-014, 3.507529e-011, 6.417138e-011,
  0, 0, 0, 0,
  1.711744e-014, 9.951233e-014, 3.273234e-011, 7.335831e-011,
  0, 0, 0, 0,
  1.623791e-014, 3.930501e-014, 3.775547e-011, 5.643411e-011,
  0, 0, 0, 0,
  1.340937e-014, 3.926611e-014, 4.518033e-011, 7.517006e-011,
  0, 0, 0, 0,
  5.847035e-014, 5.239359e-014, 6.410544e-011, 1.000722e-010,
  0, 0, 0, 0,
  3.209889e-014, 1.308194e-013, 8.194365e-011, 1.143022e-010,
  0, 0, 0, 0,
  2.993518e-014, 1.018726e-013, 1.048101e-010, 1.71462e-010,
  0, 0, 0, 0,
  3.173854e-014, 1.303098e-013, 1.837523e-010, 2.542037e-010,
  0, 0, 0, 0,
  3.656111e-014, 7.927292e-014, 1.026425e-010, 1.840256e-010,
  0, 0, 0, 0,
  6.079716e-014, 5.042669e-014, 1.461975e-010, 2.385817e-010,
  0, 0, 0, 0,
  3.212415e-014, 3.382119e-014, 2.084468e-010, 3.081387e-010,
  0, 0, 0, 0,
  2.442391e-014, 1.296112e-013, 1.219305e-010, 2.146894e-010,
  0, 0, 0, 0,
  1.567579e-014, 5.091628e-014, 1.080801e-010, 1.465784e-010,
  0, 0, 0, 0,
  2.122348e-014, 5.813907e-014, 9.341494e-011, 1.509178e-010,
  0, 0, 0, 0,
  1.915426e-014, 1.405232e-014, 5.901653e-011, 9.182806e-011,
  0, 0, 0, 0,
  1.749216e-014, 7.157901e-014, 6.569464e-011, 9.815377e-011,
  0, 0, 0, 0,
  1.809963e-014, 6.243676e-014, 6.220793e-011, 9.169814e-011,
  0, 0, 0, 0,
  7.459995e-014, 6.125704e-014, 6.449885e-011, 1.077168e-010,
  0, 0, 0, 0,
  1.665984e-014, 6.161925e-014, 3.690733e-011, 7.958353e-011,
  0, 0, 0, 0,
  1.165232e-014, 4.727982e-014, 2.859468e-011, 5.889632e-011,
  0, 0, 0, 0,
  2.213065e-014, 1.216506e-013, 4.038377e-011, 9.975201e-011,
  0, 0, 0, 0,
  7.148697e-014, 8.601593e-014, 5.466847e-011, 1.168191e-010,
  0, 0, 0, 0,
  1.93937e-014, 2.879832e-014, 4.540172e-011, 9.198009e-011,
  0, 0, 0, 0,
  1.041472e-014, 2.501531e-014, 3.72982e-011, 6.937589e-011,
  0, 0, 0, 0,
  2.784232e-014, 9.187687e-014, 9.012428e-011, 1.307148e-010,
  0, 0, 0, 0,
  2.631535e-014, 1.352473e-013, 6.628417e-011, 1.291544e-010,
  0, 0, 0, 0,
  2.939701e-014, 1.112929e-013, 7.862802e-011, 1.248822e-010,
  0, 0, 0, 0,
  3.218991e-014, 6.598022e-014, 8.730151e-011, 1.269415e-010,
  0, 0, 0, 0,
  5.211957e-014, 2.691881e-013, 1.989847e-010, 3.137045e-010,
  0, 0, 0, 0,
  3.332376e-014, 1.276518e-013, 1.822452e-010, 2.541742e-010,
  0, 0, 0, 0,
  4.454186e-014, 6.851344e-014, 1.416442e-010, 2.069997e-010,
  0, 0, 0, 0,
  5.550255e-014, 2.597016e-013, 1.932855e-010, 3.264531e-010,
  0, 0, 0, 0,
  3.342781e-014, 1.446011e-013, 2.039349e-010, 3.107247e-010,
  0, 0, 0, 0,
  3.349665e-014, 1.112551e-013, 7.470684e-011, 1.441586e-010,
  0, 0, 0, 0,
  4.717853e-015, 2.750218e-015, 2.81688e-012, 4.052502e-012,
  0, 0, 0, 0,
  2.169994e-014, 4.225446e-015, 3.455529e-011, 2.948821e-011,
  0, 0, 0, 0,
  7.330292e-014, 1.16507e-014, 5.234679e-012, 5.049589e-012,
  0, 0, 0, 0,
  6.941511e-015, 6.371537e-015, 7.051245e-012, 1.044517e-011,
  0, 0, 0, 0,
  4.781678e-015, 7.772056e-015, 4.616444e-012, 6.754258e-012,
  0, 0, 0, 0,
  3.225011e-015, 5.982376e-015, 1.028108e-011, 7.972224e-012,
  0, 0, 0, 0,
  7.895145e-014, 1.302029e-014, 7.394849e-012, 9.490972e-012,
  0, 0, 0, 0,
  5.770832e-015, 1.52764e-014, 8.779808e-012, 1.172594e-011,
  0, 0, 0, 0,
  7.801718e-014, 1.280074e-014, 1.991547e-011, 2.147945e-011,
  0, 0, 0, 0,
  8.099303e-014, 1.375859e-013, 1.851108e-011, 1.999458e-011,
  0, 0, 0, 0,
  7.419305e-014, 1.367716e-014, 3.797779e-012, 5.587271e-012,
  0, 0, 0, 0,
  9.317909e-015, 2.486794e-015, 4.167226e-012, 4.97381e-012,
  0, 0, 0, 0,
  6.7318e-015, 4.001635e-015, 5.759899e-012, 7.491809e-012,
  0, 0, 0, 0,
  1.02766e-014, 3.200344e-015, 6.094717e-012, 8.650008e-012,
  0, 0, 0, 0,
  6.587146e-015, 2.517999e-015, 5.654977e-012, 7.713778e-012,
  0, 0, 0, 0,
  1.648372e-014, 5.072086e-015, 1.053141e-011, 1.359072e-011,
  0, 0, 0, 0,
  2.004801e-014, 5.663872e-015, 1.577705e-011, 1.837622e-011,
  0, 0, 0, 0,
  3.026063e-015, 2.875147e-015, 2.919408e-012, 3.833877e-012,
  0, 0, 0, 0,
  5.173801e-015, 4.263649e-015, 4.189893e-012, 4.649094e-012,
  0, 0, 0, 0,
  8.795358e-015, 4.809097e-015, 4.012449e-012, 5.557165e-012,
  0, 0, 0, 0,
  1.271532e-014, 2.989232e-015, 9.431754e-012, 1.307213e-011,
  0, 0, 0, 0,
  1.100844e-014, 3.303671e-015, 7.059903e-012, 7.127443e-012,
  0, 0, 0, 0,
  1.560693e-014, 4.730341e-015, 6.776352e-012, 8.279262e-012,
  0, 0, 0, 0,
  6.981143e-014, 1.273284e-014, 7.008443e-012, 1.080313e-011,
  0, 0, 0, 0,
  1.074595e-014, 9.779552e-015, 5.975145e-012, 9.107163e-012,
  0, 0, 0, 0,
  5.040741e-015, 7.04699e-015, 4.077239e-012, 5.123982e-012,
  0, 0, 0, 0,
  9.969638e-015, 1.602524e-014, 4.946165e-012, 6.717646e-012,
  0, 0, 0, 0,
  8.441949e-014, 1.360433e-014, 1.326432e-011, 1.741754e-011,
  0, 0, 0, 0,
  6.821989e-015, 8.264407e-015, 6.920895e-012, 8.939152e-012,
  0, 0, 0, 0,
  1.065973e-014, 5.979703e-015, 1.041962e-011, 1.205233e-011,
  0, 0, 0, 0,
  3.705457e-015, 1.719727e-015, 2.776712e-012, 4.048189e-012,
  0, 0, 0, 0,
  6.342684e-015, 2.526469e-015, 1.187729e-011, 5.896059e-011,
  0, 0, 0, 0,
  1.304786e-014, 4.152864e-015, 8.636679e-012, 1.099976e-011,
  0, 0, 0, 0,
  1.113024e-014, 3.172598e-015, 4.416568e-012, 3.964429e-012,
  0, 0, 0, 0,
  5.417134e-015, 4.704028e-015, 1.041304e-011, 7.734429e-012,
  0, 0, 0, 0,
  5.144314e-014, 1.175725e-014, 8.679465e-012, 1.323684e-011,
  0, 0, 0, 0,
  6.373369e-014, 1.029271e-014, 7.831052e-012, 1.001941e-011,
  0, 0, 0, 0,
  6.883482e-015, 3.286887e-015, 2.899892e-012, 2.901735e-012,
  0, 0, 0, 0,
  9.186071e-015, 2.921265e-015, 2.628072e-012, 2.375967e-012,
  0, 0, 0, 0,
  1.342483e-014, 2.821858e-015, 3.515357e-012, 3.180638e-012,
  0, 0, 0, 0,
  6.650034e-014, 1.155519e-014, 4.06726e-012, 5.20589e-012,
  0, 0, 0, 0,
  1.447743e-014, 3.537263e-015, 9.002563e-012, 1.171104e-011,
  0, 0, 0, 0,
  9.92834e-015, 3.036616e-015, 6.560547e-012, 7.661964e-012,
  0, 0, 0, 0,
  6.903792e-015, 3.109175e-015, 5.352252e-012, 5.544086e-012,
  0, 0, 0, 0,
  8.403227e-014, 1.32247e-014, 2.442428e-012, 2.692112e-012,
  0, 0, 0, 0,
  3.793028e-015, 4.699201e-015, 4.577197e-012, 4.614873e-012,
  0, 0, 0, 0,
  2.461448e-015, 1.069907e-014, 5.666865e-012, 1.456585e-011,
  0, 0, 0, 0,
  5.231054e-015, 5.226579e-015, 3.490064e-012, 4.462419e-012,
  0, 0, 0, 0,
  8.991589e-014, 3.502228e-014, 8.877774e-012, 9.625838e-012,
  0, 0, 0, 0,
  1.405718e-014, 5.999192e-015, 1.227781e-011, 1.313522e-011,
  0, 0, 0, 0,
  6.793225e-015, 5.73665e-015, 3.421141e-012, 5.35519e-012,
  0, 0, 0, 0,
  3.17884e-015, 4.079331e-015, 1.837736e-012, 3.138901e-012,
  0, 0, 0, 0,
  4.398835e-014, 8.951698e-015, 2.578114e-012, 4.835008e-012,
  0, 0, 0, 0,
  3.393906e-014, 1.268944e-014, 5.734027e-012, 9.310142e-012,
  0, 0, 0, 0,
  2.966007e-015, 2.003152e-015, 2.24567e-012, 3.090799e-012,
  0, 0, 0, 0,
  6.959477e-015, 2.360591e-015, 3.683368e-012, 3.795085e-012,
  0, 0, 0, 0,
  2.3648e-014, 5.47648e-015, 4.680381e-012, 5.715521e-012,
  0, 0, 0, 0,
  6.082186e-014, 1.050374e-014, 6.036958e-012, 8.398031e-012,
  0, 0, 0, 0,
  6.513997e-015, 4.591763e-015, 3.600457e-012, 3.598901e-012,
  0, 0, 0, 0,
  3.126923e-015, 2.060524e-015, 2.021821e-012, 2.291461e-012,
  0, 0, 0, 0,
  2.655934e-015, 4.092173e-015, 2.493609e-012, 3.001514e-012,
  0, 0, 0, 0,
  2.266697e-015, 2.23642e-015, 2.191133e-012, 2.809541e-012,
  0, 0, 0, 0,
  4.010466e-015, 1.97059e-015, 2.032058e-012, 3.373834e-012,
  0, 0, 0, 0,
  2.404577e-015, 1.904929e-015, 2.762136e-012, 2.760745e-012,
  0, 0, 0, 0,
  2.128259e-015, 3.290851e-015, 2.165558e-012, 1.945193e-012,
  0, 0, 0, 0,
  8.908613e-014, 1.614873e-014, 2.978678e-012, 5.998772e-012,
  0, 0, 0, 0,
  3.77482e-015, 5.301117e-015, 2.322003e-012, 3.673873e-012,
  0, 0, 0, 0,
  5.249906e-015, 1.341496e-014, 1.431642e-011, 2.047164e-011,
  0, 0, 0, 0,
  1.026404e-014, 1.263009e-014, 1.424826e-011, 2.129256e-011,
  0, 0, 0, 0,
  6.088352e-014, 1.01694e-014, 9.995398e-012, 9.239652e-012,
  0, 0, 0, 0,
  1.775382e-014, 4.903256e-015, 3.205651e-012, 3.481131e-012,
  0, 0, 0, 0,
  6.286717e-015, 5.14457e-015, 1.065365e-011, 1.225663e-011,
  0, 0, 0, 0,
  6.030909e-015, 3.673516e-015, 4.109702e-012, 5.043456e-012,
  0, 0, 0, 0,
  3.506923e-014, 6.886153e-015, 3.213273e-012, 3.82886e-012,
  0, 0, 0, 0,
  5.051115e-014, 8.112409e-015, 3.438097e-012, 3.128216e-012,
  0, 0, 0, 0,
  2.863118e-015, 3.299838e-015, 3.544973e-012, 3.697382e-012,
  0, 0, 0, 0,
  5.192993e-015, 4.461317e-015, 3.031427e-012, 2.586276e-012,
  0, 0, 0, 0,
  5.78092e-015, 4.144372e-015, 3.747098e-012, 6.556462e-012,
  0, 0, 0, 0,
  8.472297e-015, 1.290463e-014, 6.927315e-012, 1.043207e-011,
  0, 0, 0, 0,
  6.67248e-015, 7.026946e-015, 5.458167e-012, 6.469076e-012,
  0, 0, 0, 0,
  1.218484e-014, 9.622728e-015, 1.260997e-011, 1.543525e-011,
  0, 0, 0, 0,
  1.835712e-014, 1.073049e-014, 1.007562e-011, 1.635907e-011,
  0, 0, 0, 0,
  9.217175e-014, 1.861478e-014, 6.978967e-012, 1.047673e-011,
  0, 0, 0, 0,
  1.017285e-014, 1.946966e-014, 1.293126e-011, 2.174379e-011,
  0, 0, 0, 0,
  8.958305e-015, 1.599511e-014, 7.836298e-012, 1.213151e-011,
  0, 0, 0, 0,
  9.046463e-015, 9.495399e-015, 7.305308e-012, 7.690637e-012,
  0, 0, 0, 0,
  7.527988e-014, 1.431885e-014, 6.547824e-012, 8.219167e-012,
  0, 0, 0, 0,
  1.332547e-014, 8.564719e-015, 6.870566e-012, 7.542686e-012,
  0, 0, 0, 0,
  7.107785e-015, 8.488133e-015, 7.409053e-012, 1.021687e-011,
  0, 0, 0, 0,
  9.439829e-015, 1.571104e-014, 9.043786e-012, 1.523687e-011,
  0, 0, 0, 0,
  5.311934e-014, 1.845531e-014, 6.146366e-012, 1.120561e-011,
  0, 0, 0, 0,
  3.313521e-014, 1.452217e-014, 5.229723e-012, 9.863927e-012,
  0, 0, 0, 0,
  6.894951e-015, 1.446003e-014, 7.362303e-012, 1.602989e-011,
  0, 0, 0, 0,
  7.7982e-015, 8.504871e-015, 1.221526e-011, 1.504983e-011,
  0, 0, 0, 0,
  1.034759e-014, 1.007645e-014, 3.485405e-012, 6.371562e-012,
  0, 0, 0, 0,
  9.205856e-015, 8.065349e-015, 4.795079e-012, 8.004109e-012,
  0, 0, 0, 0,
  1.062811e-014, 4.278039e-015, 4.457481e-012, 5.45959e-012,
  0, 0, 0, 0,
  5.748644e-015, 5.944782e-015, 6.364591e-012, 6.89719e-012,
  0, 0, 0, 0,
  4.095985e-015, 7.863922e-015, 8.123313e-012, 8.628227e-012,
  0, 0, 0, 0,
  3.820981e-015, 7.34768e-015, 4.495807e-012, 5.716565e-012,
  0, 0, 0, 0,
  2.298869e-015, 3.278555e-015, 2.61005e-012, 2.872963e-012,
  0, 0, 0, 0,
  4.05369e-015, 9.926911e-015, 3.327445e-012, 2.866119e-012,
  0, 0, 0, 0,
  2.519858e-013, 3.938366e-014, 4.618735e-011, 6.174655e-011,
  0, 0, 0, 0,
  6.008245e-014, 1.114718e-014, 6.036355e-011, 6.704001e-011,
  0, 0, 0, 0,
  2.072501e-014, 1.415147e-014, 3.288763e-011, 4.507607e-011,
  0, 0, 0, 0,
  1.01644e-013, 3.174675e-014, 7.535189e-011, 1.173963e-010,
  0, 0, 0, 0,
  7.355618e-015, 8.568125e-015, 4.895536e-012, 9.000848e-012,
  0, 0, 0, 0,
  1.374811e-014, 9.364886e-015, 6.719942e-012, 8.843292e-012,
  0, 0, 0, 0,
  1.767421e-014, 9.32148e-015, 2.082726e-011, 2.620343e-011,
  0, 0, 0, 0,
  2.172284e-014, 1.151997e-014, 5.204863e-012, 1.148871e-011,
  0, 0, 0, 0,
  1.4145e-014, 1.069368e-014, 5.552336e-012, 1.056667e-011,
  0, 0, 0, 0,
  1.893561e-014, 8.538682e-015, 4.610862e-012, 8.311193e-012,
  0, 0, 0, 0,
  1.888721e-014, 8.011033e-015, 3.922595e-012, 6.105047e-012,
  0, 0, 0, 0,
  4.88133e-014, 1.128888e-014, 5.060845e-012, 1.263137e-011,
  0, 0, 0, 0,
  5.943447e-014, 1.429535e-014, 1.658472e-011, 1.887013e-011,
  0, 0, 0, 0,
  1.067336e-013, 1.998649e-014, 1.586937e-011, 1.820128e-011,
  0, 0, 0, 0,
  5.380883e-014, 1.563876e-014, 4.595116e-012, 9.430111e-012,
  0, 0, 0, 0,
  8.228373e-014, 2.726168e-014, 5.98192e-012, 1.283516e-011,
  0, 0, 0, 0,
  1.614639e-013, 3.710656e-014, 7.278852e-012, 1.969608e-011,
  0, 0, 0, 0,
  5.659047e-013, 9.382095e-014, 1.089434e-011, 5.037367e-011,
  0, 0, 0, 0,
  2.699597e-013, 6.252652e-014, 9.252871e-012, 3.077141e-011,
  0, 0, 0, 0,
  5.158206e-013, 9.958095e-014, 1.68701e-011, 6.869372e-011,
  0, 0, 0, 0,
  6.605884e-013, 1.403306e-013, 2.100539e-011, 9.232535e-011,
  0, 0, 0, 0,
  1.381007e-012, 2.912341e-013, 4.111235e-011, 1.898145e-010,
  0, 0, 0, 0,
  2.130403e-012, 4.436273e-013, 1.186611e-010, 4.451213e-010,
  0, 0, 0, 0,
  2.361569e-012, 5.491152e-013, 9.539045e-011, 3.895418e-010,
  0, 0, 0, 0,
  4.039402e-012, 1.096833e-012, 1.898201e-010, 7.475596e-010,
  0, 0, 0, 0,
  7.038811e-012, 2.286916e-012, 6.742611e-010, 1.709829e-009,
  0, 0, 0, 0,
  1.397733e-011, 4.30255e-012, 1.437062e-009, 7.299715e-009,
  0, 0, 0, 0,
  1.744823e-011, 4.868949e-012, 1.088757e-009, 3.844548e-009,
  0, 0, 0, 0,
  8.795401e-012, 3.519726e-012, 8.209537e-010, 2.51012e-009,
  0, 0, 0, 0,
  1.312297e-011, 3.708503e-012, 8.522967e-010, 2.938463e-009,
  0, 0, 0, 0,
  1.346471e-011, 5.079367e-012, 1.002368e-009, 3.762032e-009,
  0, 0, 0, 0,
  4.479325e-012, 2.341829e-012, 3.710635e-010, 1.522317e-009,
  0, 0, 0, 0,
  3.040786e-012, 6.712982e-013, 1.285801e-010, 5.479052e-010,
  0, 0, 0, 0,
  1.81563e-012, 4.827384e-013, 6.631586e-011, 2.866074e-010,
  0, 0, 0, 0,
  1.696539e-012, 4.721876e-013, 5.548245e-011, 2.606157e-010,
  0, 0, 0, 0,
  1.092297e-012, 3.452843e-013, 3.444619e-011, 1.622303e-010,
  0, 0, 0, 0,
  7.240118e-013, 1.874751e-013, 3.031086e-011, 9.69952e-011,
  0, 0, 0, 0,
  3.322709e-013, 1.928981e-013, 2.15472e-011, 3.82218e-011,
  0, 0, 0, 0,
  3.828948e-013, 2.484846e-013, 2.192707e-011, 6.480069e-011,
  0, 0, 0, 0,
  3.06737e-013, 1.26275e-013, 2.083861e-011, 8.753248e-011,
  0, 0, 0, 0,
  2.435325e-013, 4.926596e-014, 7.896289e-012, 2.49812e-011,
  0, 0, 0, 0,
  8.81977e-014, 4.136943e-014, 1.003191e-011, 2.606555e-011,
  0, 0, 0, 0,
  1.239416e-013, 3.993009e-014, 1.118461e-011, 2.634097e-011,
  0, 0, 0, 0,
  8.086973e-014, 2.295658e-013, 4.556213e-011, 1.286582e-010,
  0, 0, 0, 0,
  3.688697e-014, 1.734733e-014, 5.377311e-012, 1.192115e-011,
  0, 0, 0, 0,
  3.331639e-014, 1.539507e-014, 9.396354e-012, 1.455176e-011,
  0, 0, 0, 0,
  2.268868e-014, 2.158882e-014, 9.473854e-012, 1.824384e-011,
  0, 0, 0, 0,
  3.805972e-014, 3.57039e-014, 1.342803e-011, 2.511129e-011,
  0, 0, 0, 0,
  4.2122e-014, 1.398721e-013, 3.524998e-011, 9.058972e-011,
  0, 0, 0, 0,
  3.538163e-014, 1.140662e-013, 2.653699e-011, 7.265604e-011,
  0, 0, 0, 0,
  6.37613e-014, 3.908904e-013, 6.575157e-011, 2.212041e-010,
  0, 0, 0, 0,
  8.144281e-014, 1.394486e-013, 2.576665e-011, 8.014807e-011,
  0, 0, 0, 0,
  3.586288e-014, 1.389923e-013, 2.983478e-011, 8.648875e-011,
  0, 0, 0, 0,
  1.868591e-014, 5.092475e-014, 2.03866e-011, 3.716947e-011,
  0, 0, 0, 0,
  1.444525e-014, 4.189671e-014, 1.583607e-011, 3.204744e-011,
  0, 0, 0, 0,
  1.432272e-014, 7.325928e-014, 1.981096e-011, 4.339819e-011,
  0, 0, 0, 0,
  1.317384e-014, 2.968646e-014, 9.86273e-012, 1.997355e-011,
  0, 0, 0, 0,
  7.819081e-015, 1.328137e-014, 1.342698e-011, 1.475493e-011,
  0, 0, 0, 0,
  9.245536e-015, 1.193838e-014, 7.503216e-012, 1.071618e-011,
  0, 0, 0, 0,
  1.098748e-014, 5.773424e-014, 1.776506e-011, 4.404856e-011,
  0, 0, 0, 0,
  1.11625e-014, 2.067659e-014, 8.924456e-012, 1.758987e-011,
  0, 0, 0, 0,
  1.14156e-014, 2.092798e-014, 7.042083e-012, 1.570304e-011,
  0, 0, 0, 0,
  6.994077e-015, 2.351618e-014, 9.03574e-012, 1.561463e-011,
  0, 0, 0, 0,
  9.735097e-014, 2.744072e-014, 1.805647e-011, 2.359532e-011,
  0, 0, 0, 0,
  1.148864e-014, 5.867104e-014, 1.359492e-011, 3.741719e-011,
  0, 0, 0, 0,
  2.971889e-014, 7.323685e-014, 2.406035e-011, 3.895984e-011,
  0, 0, 0, 0,
  2.863757e-014, 1.314371e-013, 2.900234e-011, 6.842471e-011,
  0, 0, 0, 0,
  5.375073e-014, 3.398193e-013, 5.497317e-011, 1.630496e-010,
  0, 0, 0, 0,
  9.896266e-014, 2.993236e-013, 7.025183e-011, 1.797111e-010,
  0, 0, 0, 0,
  4.19682e-014, 2.354576e-013, 7.087712e-011, 1.810999e-010,
  0, 0, 0, 0,
  5.164445e-014, 2.978181e-013, 5.661034e-011, 1.735543e-010,
  0, 0, 0, 0,
  2.195828e-014, 1.049497e-013, 2.029809e-011, 5.306024e-011,
  0, 0, 0, 0,
  6.673326e-014, 1.01507e-013, 3.167717e-011, 7.522904e-011,
  0, 0, 0, 0,
  1.616686e-014, 3.630918e-014, 1.796056e-011, 3.263792e-011,
  0, 0, 0, 0,
  7.109419e-015, 2.136208e-014, 1.143812e-011, 1.952058e-011,
  0, 0, 0, 0,
  1.663378e-014, 9.842844e-014, 2.010865e-011, 6.075988e-011,
  0, 0, 0, 0,
  5.705638e-014, 1.805136e-013, 2.460595e-011, 8.797265e-011,
  0, 0, 0, 0,
  3.446757e-014, 5.628811e-014, 1.184044e-011, 2.866958e-011,
  0, 0, 0, 0,
  2.946136e-014, 1.127641e-013, 2.705681e-011, 7.221371e-011,
  0, 0, 0, 0,
  3.005133e-014, 1.031494e-013, 2.113604e-011, 5.877097e-011,
  0, 0, 0, 0,
  6.284934e-014, 3.944222e-013, 6.733748e-011, 2.104746e-010,
  0, 0, 0, 0,
  2.037138e-014, 8.057992e-014, 3.832761e-011, 7.967248e-011,
  0, 0, 0, 0,
  6.442137e-014, 4.05153e-013, 6.164275e-011, 1.903297e-010,
  0, 0, 0, 0,
  3.464892e-014, 1.769433e-013, 3.89587e-011, 1.064057e-010,
  0, 0, 0, 0,
  6.983925e-014, 4.337851e-013, 9.573678e-011, 2.762365e-010,
  0, 0, 0, 0,
  1.016498e-013, 1.748241e-013, 3.821624e-011, 1.015338e-010,
  0, 0, 0, 0,
  3.955594e-014, 2.084321e-013, 7.115062e-011, 1.735733e-010,
  0, 0, 0, 0,
  4.546246e-014, 1.515756e-013, 4.686644e-011, 1.080443e-010,
  0, 0, 0, 0,
  4.356008e-014, 2.720395e-013, 4.785632e-011, 1.46808e-010,
  0, 0, 0, 0,
  7.102065e-014, 6.858429e-014, 1.23926e-011, 3.37574e-011,
  0, 0, 0, 0,
  1.284964e-014, 3.3624e-014, 1.445538e-011, 2.388288e-011,
  0, 0, 0, 0,
  1.034121e-014, 2.594951e-014, 2.241317e-011, 3.728267e-011,
  0, 0, 0, 0,
  9.416764e-015, 4.506752e-014, 1.456586e-011, 2.884129e-011,
  0, 0, 0, 0,
  5.97694e-014, 2.149767e-014, 9.310068e-012, 1.705019e-011,
  0, 0, 0, 0,
  2.172831e-014, 1.517743e-014, 8.203362e-012, 1.20261e-011,
  0, 0, 0, 0,
  1.177876e-014, 2.42808e-014, 8.27842e-012, 1.409102e-011,
  0, 0, 0, 0,
  5.322282e-015, 2.509576e-014, 6.438214e-012, 1.341752e-011,
  0, 0, 0, 0,
  7.140234e-015, 2.300832e-014, 8.967646e-012, 1.588015e-011,
  0, 0, 0, 0,
  8.937774e-015, 3.734629e-014, 1.459617e-011, 2.517343e-011,
  0, 0, 0, 0,
  9.322235e-015, 2.204197e-014, 1.031567e-011, 1.883644e-011,
  0, 0, 0, 0,
  1.265671e-014, 2.08331e-014, 9.904177e-012, 1.721182e-011,
  0, 0, 0, 0,
  3.976172e-014, 2.283416e-013, 3.392061e-011, 1.038397e-010,
  0, 0, 0, 0,
  1.220095e-013, 3.57138e-013, 5.199511e-011, 1.515133e-010,
  0, 0, 0, 0,
  4.775803e-014, 2.817187e-013, 4.569306e-011, 1.364165e-010,
  0, 0, 0, 0,
  8.594736e-014, 5.401633e-013, 9.197154e-011, 2.638589e-010,
  0, 0, 0, 0,
  7.563625e-014, 4.196079e-013, 8.591327e-011, 1.91663e-010,
  0, 0, 0, 0,
  1.015353e-013, 4.704246e-013, 8.042582e-011, 2.492782e-010,
  0, 0, 0, 0,
  9.467882e-014, 4.875124e-013, 8.999923e-011, 2.05163e-010,
  0, 0, 0, 0,
  1.594636e-013, 9.463206e-013, 2.099938e-010, 5.496082e-010,
  0, 0, 0, 0,
  7.729397e-014, 3.851767e-013, 8.246542e-011, 1.706167e-010,
  0, 0, 0, 0,
  9.553333e-014, 3.592146e-013, 1.170155e-010, 2.700583e-010,
  0, 0, 0, 0,
  6.627173e-014, 2.312605e-013, 1.055583e-010, 2.226831e-010,
  0, 0, 0, 0,
  9.327904e-014, 3.199122e-013, 1.532874e-010, 2.917308e-010,
  0, 0, 0, 0,
  6.730781e-014, 1.390276e-013, 1.357788e-010, 2.397323e-010,
  0, 0, 0, 0,
  1.124202e-013, 3.555018e-013, 2.710605e-010, 4.278082e-010,
  0, 0, 0, 0,
  9.034433e-014, 2.532541e-013, 1.356781e-010, 2.266503e-010,
  0, 0, 0, 0,
  1.594692e-013, 7.315274e-013, 1.811039e-010, 4.838694e-010,
  0, 0, 0, 0,
  8.544559e-014, 2.807979e-013, 1.224617e-010, 2.482015e-010,
  0, 0, 0, 0,
  4.174342e-014, 1.314162e-013, 7.688707e-011, 1.381482e-010,
  0, 0, 0, 0,
  6.335978e-014, 1.642557e-013, 4.965329e-011, 9.695943e-011,
  0, 0, 0, 0,
  4.208602e-014, 1.025617e-013, 8.827306e-011, 1.247319e-010,
  0, 0, 0, 0,
  4.124046e-014, 6.07212e-014, 4.732825e-011, 7.201674e-011,
  0, 0, 0, 0,
  2.710876e-014, 1.887223e-014, 2.101689e-011, 3.404512e-011,
  0, 0, 0, 0,
  8.46345e-014, 2.533885e-014, 3.860474e-011, 4.965149e-011,
  0, 0, 0, 0,
  2.160288e-014, 2.144624e-014, 1.271697e-011, 1.71298e-011,
  0, 0, 0, 0,
  1.490179e-014, 1.024344e-014, 7.419219e-012, 1.250271e-011,
  0, 0, 0, 0,
  1.534506e-014, 9.440312e-015, 9.672587e-012, 1.527388e-011,
  0, 0, 0, 0,
  1.650529e-014, 8.980109e-015, 6.96464e-012, 1.117646e-011,
  0, 0, 0, 0,
  1.284323e-014, 9.596873e-015, 8.597914e-012, 1.347948e-011,
  0, 0, 0, 0,
  1.297992e-014, 1.150705e-014, 7.963237e-012, 1.079776e-011,
  0, 0, 0, 0,
  2.068092e-014, 2.130207e-014, 8.092255e-012, 1.551283e-011,
  0, 0, 0, 0,
  4.735901e-014, 2.252389e-014, 1.029687e-011, 1.876161e-011,
  0, 0, 0, 0,
  2.900093e-014, 8.379019e-014, 1.475107e-011, 4.057403e-011,
  0, 0, 0, 0,
  4.526848e-014, 8.551013e-014, 2.435728e-011, 5.82942e-011,
  0, 0, 0, 0,
  1.808962e-014, 2.530812e-014, 2.328132e-011, 3.158621e-011,
  0, 0, 0, 0,
  3.568623e-014, 1.570235e-014, 1.568583e-011, 2.462463e-011,
  0, 0, 0, 0,
  6.41449e-014, 3.041115e-014, 2.328492e-011, 3.501124e-011,
  0, 0, 0, 0,
  4.774367e-014, 4.86476e-014, 4.694967e-011, 7.869904e-011,
  0, 0, 0, 0,
  3.85654e-014, 1.699307e-014, 6.513051e-011, 1.090531e-010,
  0, 0, 0, 0,
  5.425204e-014, 3.00278e-014, 8.932591e-011, 1.499663e-010,
  0, 0, 0, 0,
  4.97806e-014, 2.836079e-014, 1.372332e-010, 1.781791e-010,
  0, 0, 0, 0,
  3.169405e-014, 2.729709e-014, 7.262432e-011, 1.056701e-010,
  0, 0, 0, 0,
  5.440788e-014, 2.167432e-014, 9.543193e-011, 1.583439e-010,
  0, 0, 0, 0,
  9.255898e-014, 3.991008e-014, 1.383081e-010, 2.240018e-010,
  0, 0, 0, 0,
  9.747929e-014, 4.101869e-014, 1.113833e-010, 1.994816e-010,
  0, 0, 0, 0,
  7.132572e-014, 3.527116e-014, 1.434247e-010, 2.541856e-010,
  0, 0, 0, 0,
  1.344189e-013, 6.396508e-014, 2.241814e-010, 4.252561e-010,
  0, 0, 0, 0,
  1.033007e-013, 1.893728e-013, 1.986552e-010, 3.874904e-010,
  0, 0, 0, 0,
  1.177609e-013, 2.587338e-013, 4.565572e-010, 7.512755e-010,
  0, 0, 0, 0,
  1.169808e-013, 6.212771e-013, 1.341113e-010, 3.070678e-010,
  0, 0, 0, 0,
  9.457433e-014, 3.555526e-013, 1.758019e-010, 3.546786e-010,
  0, 0, 0, 0,
  8.367614e-014, 3.43255e-013, 2.969293e-010, 4.240573e-010,
  0, 0, 0, 0,
  1.008334e-013, 3.898854e-013, 3.136273e-010, 5.65706e-010,
  0, 0, 0, 0,
  7.609724e-014, 7.399874e-014, 1.576154e-010, 2.609286e-010,
  0, 0, 0, 0,
  5.762695e-014, 2.030122e-013, 5.991948e-011, 1.29557e-010,
  0, 0, 0, 0,
  3.606089e-014, 6.669579e-014, 3.357964e-011, 5.524486e-011,
  0, 0, 0, 0,
  8.52987e-014, 5.555642e-014, 1.370871e-010, 2.131386e-010,
  0, 0, 0, 0,
  6.52669e-014, 2.501012e-014, 1.689672e-011, 2.556335e-011,
  0, 0, 0, 0,
  3.797302e-014, 3.024339e-014, 6.37936e-011, 1.057072e-010,
  0, 0, 0, 0,
  1.556298e-014, 2.701851e-014, 2.212989e-011, 3.44022e-011,
  0, 0, 0, 0,
  3.206537e-014, 2.089371e-014, 4.227595e-011, 6.547343e-011,
  0, 0, 0, 0,
  6.241238e-014, 3.4232e-014, 3.38413e-011, 5.430078e-011,
  0, 0, 0, 0,
  2.81166e-014, 3.556896e-014, 3.28545e-011, 4.798655e-011,
  0, 0, 0, 0,
  3.113757e-014, 1.037063e-013, 7.119694e-011, 1.052409e-010,
  0, 0, 0, 0,
  1.061665e-013, 6.172685e-013, 9.368056e-011, 2.645679e-010,
  0, 0, 0, 0,
  3.788665e-014, 5.690026e-014, 5.408915e-011, 9.893794e-011,
  0, 0, 0, 0,
  4.119166e-014, 7.842261e-014, 6.320277e-011, 1.103429e-010,
  0, 0, 0, 0,
  7.663251e-014, 3.938968e-013, 7.421731e-011, 2.077571e-010,
  0, 0, 0, 0,
  7.322951e-014, 3.627529e-013, 9.372284e-011, 2.140403e-010,
  0, 0, 0, 0,
  7.29113e-014, 1.674483e-013, 9.928466e-011, 1.754962e-010,
  0, 0, 0, 0,
  5.26934e-014, 1.793451e-013, 8.421697e-011, 1.647082e-010,
  0, 0, 0, 0,
  2.944444e-014, 9.423731e-014, 4.861124e-011, 6.510746e-011,
  0, 0, 0, 0,
  2.839252e-014, 8.041454e-014, 4.359888e-011, 8.867131e-011,
  0, 0, 0, 0,
  6.934438e-014, 1.267992e-013, 7.462905e-011, 1.321629e-010,
  0, 0, 0, 0,
  5.759147e-014, 1.799996e-013, 2.444824e-010, 2.856111e-010,
  0, 0, 0, 0,
  4.341133e-014, 1.448166e-013, 5.831871e-011, 1.059146e-010,
  0, 0, 0, 0,
  4.920602e-014, 1.141741e-013, 7.039958e-011, 1.067002e-010,
  0, 0, 0, 0,
  7.109827e-014, 1.422828e-013, 1.185701e-010, 1.862143e-010,
  0, 0, 0, 0,
  8.396128e-014, 4.051771e-014, 2.648235e-011, 4.766323e-011,
  0, 0, 0, 0,
  3.635388e-014, 8.741963e-014, 6.361346e-011, 9.395301e-011,
  0, 0, 0, 0,
  3.213914e-014, 1.725493e-013, 3.687659e-011, 9.197217e-011,
  0, 0, 0, 0,
  3.104018e-014, 1.365574e-013, 6.044786e-011, 1.020784e-010,
  0, 0, 0, 0,
  4.143556e-014, 2.234256e-013, 6.503004e-011, 1.270672e-010,
  0, 0, 0, 0,
  3.155988e-014, 1.304403e-013, 3.765869e-011, 7.264644e-011,
  0, 0, 0, 0,
  2.632081e-014, 5.260617e-014, 6.129851e-011, 9.024231e-011,
  0, 0, 0, 0,
  2.403279e-014, 6.437224e-014, 5.473401e-011, 8.953888e-011,
  0, 0, 0, 0,
  6.428809e-014, 1.105375e-013, 7.382314e-011, 1.368691e-010,
  0, 0, 0, 0,
  5.109899e-014, 1.407823e-013, 1.454143e-010, 2.149072e-010,
  0, 0, 0, 0,
  7.062675e-014, 1.620285e-013, 4.354737e-010, 6.35534e-010,
  0, 0, 0, 0,
  1.072659e-013, 1.375238e-013, 3.43972e-010, 5.734984e-010,
  0, 0, 0, 0,
  8.999575e-014, 2.637938e-013, 1.449486e-010, 2.66211e-010,
  0, 0, 0, 0,
  1.045719e-013, 7.89253e-014, 2.946506e-010, 4.730041e-010,
  0, 0, 0, 0,
  1.615995e-013, 7.030155e-014, 3.586784e-010, 6.218837e-010,
  0, 0, 0, 0,
  1.071841e-013, 2.908411e-013, 2.535792e-010, 3.974255e-010,
  0, 0, 0, 0,
  1.050245e-013, 8.851693e-014, 2.850302e-010, 4.152974e-010,
  0, 0, 0, 0,
  4.125261e-014, 8.306935e-014, 1.052569e-010, 1.423404e-010,
  0, 0, 0, 0,
  4.29866e-014, 5.50108e-014, 1.004774e-010, 1.604107e-010,
  0, 0, 0, 0,
  5.201768e-014, 8.900241e-014, 9.757578e-011, 1.322748e-010,
  0, 0, 0, 0,
  9.178877e-014, 9.485778e-014, 2.320733e-010, 3.552595e-010,
  0, 0, 0, 0,
  6.466791e-014, 6.917207e-014, 1.04534e-010, 1.489958e-010,
  0, 0, 0, 0,
  4.74153e-014, 9.941632e-014, 6.784227e-011, 1.289078e-010,
  0, 0, 0, 0,
  7.914962e-014, 1.506078e-013, 9.565383e-011, 1.831914e-010,
  0, 0, 0, 0,
  4.767047e-014, 2.304115e-013, 6.857553e-011, 1.462524e-010,
  0, 0, 0, 0,
  7.645933e-014, 5.80996e-014, 7.50374e-011, 1.32708e-010,
  0, 0, 0, 0,
  5.036995e-014, 3.549316e-014, 1.083383e-010, 1.806459e-010,
  0, 0, 0, 0,
  3.841941e-014, 6.234196e-014, 7.676002e-011, 1.264882e-010,
  0, 0, 0, 0,
  4.274576e-014, 2.044448e-013, 1.249901e-010, 2.243583e-010,
  0, 0, 0, 0,
  4.234001e-014, 1.383351e-013, 9.924114e-011, 1.840479e-010,
  0, 0, 0, 0,
  4.252316e-014, 1.118659e-013, 1.252954e-010, 2.120816e-010,
  0, 0, 0, 0,
  8.302598e-014, 1.134858e-013, 2.024864e-010, 3.184689e-010,
  0, 0, 0, 0,
  1.250611e-013, 4.79338e-013, 3.003538e-010, 5.674521e-010,
  0, 0, 0, 0,
  1.47255e-013, 1.038402e-013, 2.963278e-010, 5.431032e-010,
  0, 0, 0, 0,
  1.361629e-013, 2.189334e-013, 3.373823e-010, 6.002933e-010,
  0, 0, 0, 0,
  1.737167e-013, 3.657676e-013, 5.243133e-010, 7.518033e-010,
  0, 0, 0, 0,
  1.497879e-013, 2.973828e-013, 3.508874e-010, 6.533115e-010,
  0, 0, 0, 0,
  1.120111e-013, 2.12426e-013, 3.49869e-010, 6.26338e-010,
  0, 0, 0, 0,
  6.385969e-015, 4.23288e-015, 3.3689e-012, 4.834117e-012,
  0, 0, 0, 0,
  2.508465e-014, 4.742647e-015, 3.529406e-011, 3.019243e-011,
  0, 0, 0, 0,
  8.283883e-014, 1.33131e-014, 6.692772e-012, 7.220069e-012,
  0, 0, 0, 0,
  1.204158e-014, 1.364133e-014, 6.423606e-012, 1.132642e-011,
  0, 0, 0, 0,
  5.309931e-015, 5.670248e-015, 6.262393e-012, 6.944716e-012,
  0, 0, 0, 0,
  6.653013e-015, 6.003376e-015, 1.279321e-011, 1.896315e-011,
  0, 0, 0, 0,
  7.949199e-014, 1.429388e-014, 7.049001e-012, 1.166307e-011,
  0, 0, 0, 0,
  5.543034e-015, 1.888169e-014, 7.726219e-012, 1.525337e-011,
  0, 0, 0, 0,
  6.162996e-014, 1.035997e-014, 2.346064e-011, 4.090647e-011,
  0, 0, 0, 0,
  5.578579e-014, 1.203953e-013, 2.080995e-011, 3.676837e-011,
  0, 0, 0, 0,
  7.890141e-014, 1.919055e-014, 3.708075e-012, 4.973619e-012,
  0, 0, 0, 0,
  1.000269e-014, 3.172606e-015, 3.751606e-012, 5.323877e-012,
  0, 0, 0, 0,
  9.054963e-015, 5.789723e-015, 9.663101e-012, 1.149637e-011,
  0, 0, 0, 0,
  1.139257e-014, 2.591885e-015, 7.521326e-012, 1.010353e-011,
  0, 0, 0, 0,
  6.082201e-015, 2.511699e-015, 7.317818e-012, 1.026986e-011,
  0, 0, 0, 0,
  8.946267e-015, 4.07195e-015, 5.476717e-012, 9.856381e-012,
  0, 0, 0, 0,
  2.071177e-014, 6.073812e-015, 1.609586e-011, 2.475278e-011,
  0, 0, 0, 0,
  4.063413e-015, 3.340963e-015, 3.896823e-012, 5.724762e-012,
  0, 0, 0, 0,
  4.918417e-015, 8.150693e-015, 7.306734e-012, 1.012396e-011,
  0, 0, 0, 0,
  7.950755e-015, 4.517335e-015, 6.232732e-012, 9.098801e-012,
  0, 0, 0, 0,
  1.964669e-014, 4.700406e-015, 1.134586e-011, 1.696809e-011,
  0, 0, 0, 0,
  1.254013e-014, 3.259095e-015, 7.660842e-012, 8.536079e-012,
  0, 0, 0, 0,
  3.512263e-014, 7.847095e-015, 1.14258e-011, 1.946028e-011,
  0, 0, 0, 0,
  7.787887e-014, 1.520932e-014, 1.795532e-011, 2.832658e-011,
  0, 0, 0, 0,
  9.546959e-015, 8.220871e-015, 9.602386e-012, 1.343046e-011,
  0, 0, 0, 0,
  5.846786e-015, 5.956328e-015, 6.250004e-012, 8.81157e-012,
  0, 0, 0, 0,
  1.333431e-014, 1.1984e-014, 5.298286e-012, 7.957432e-012,
  0, 0, 0, 0,
  8.706808e-014, 1.386965e-014, 2.163607e-011, 3.808846e-011,
  0, 0, 0, 0,
  8.739675e-015, 1.033787e-014, 5.28305e-012, 8.312302e-012,
  0, 0, 0, 0,
  1.155031e-014, 6.325992e-015, 1.014254e-011, 1.339515e-011,
  0, 0, 0, 0,
  2.877507e-015, 2.510213e-015, 3.98147e-012, 4.354237e-012,
  0, 0, 0, 0,
  2.089004e-014, 5.487653e-015, 1.106225e-011, 4.761886e-011,
  0, 0, 0, 0,
  1.2477e-014, 4.138545e-015, 7.963574e-012, 1.381693e-011,
  0, 0, 0, 0,
  2.013071e-014, 4.261902e-015, 6.70679e-012, 1.277834e-011,
  0, 0, 0, 0,
  1.273583e-014, 7.479616e-015, 7.985961e-012, 1.272432e-011,
  0, 0, 0, 0,
  5.197769e-014, 1.834046e-014, 9.855103e-012, 1.547189e-011,
  0, 0, 0, 0,
  6.341251e-014, 1.153513e-014, 1.432734e-011, 2.327352e-011,
  0, 0, 0, 0,
  7.701313e-015, 2.593699e-015, 3.618637e-012, 6.690732e-012,
  0, 0, 0, 0,
  8.767573e-015, 3.003534e-015, 2.651744e-012, 3.845091e-012,
  0, 0, 0, 0,
  1.359302e-014, 3.117951e-015, 2.496749e-012, 3.425382e-012,
  0, 0, 0, 0,
  7.044374e-014, 1.232316e-014, 4.439289e-012, 6.788688e-012,
  0, 0, 0, 0,
  2.216626e-014, 4.506093e-015, 4.481557e-012, 5.403443e-012,
  0, 0, 0, 0,
  1.113324e-014, 3.428886e-015, 4.683119e-012, 6.814261e-012,
  0, 0, 0, 0,
  7.100463e-015, 3.937477e-015, 4.60362e-012, 6.359295e-012,
  0, 0, 0, 0,
  8.765082e-014, 1.416918e-014, 2.989002e-012, 3.207091e-012,
  0, 0, 0, 0,
  6.947604e-015, 1.075611e-014, 3.25715e-012, 5.6257e-012,
  0, 0, 0, 0,
  5.866698e-015, 2.476581e-014, 6.029642e-012, 1.23279e-011,
  0, 0, 0, 0,
  4.321664e-015, 6.48851e-015, 4.14563e-012, 5.960952e-012,
  0, 0, 0, 0,
  1.027911e-013, 2.161949e-014, 1.108696e-011, 1.799939e-011,
  0, 0, 0, 0,
  1.670105e-014, 5.408344e-015, 1.770865e-011, 2.14025e-011,
  0, 0, 0, 0,
  6.878122e-015, 9.574759e-015, 4.959653e-012, 8.46171e-012,
  0, 0, 0, 0,
  2.986269e-015, 5.633179e-015, 2.147884e-012, 2.452931e-012,
  0, 0, 0, 0,
  4.6385e-014, 1.110052e-014, 2.629025e-012, 4.616185e-012,
  0, 0, 0, 0,
  3.584703e-014, 9.806168e-015, 2.797713e-012, 5.535693e-012,
  0, 0, 0, 0,
  2.555385e-015, 3.051576e-015, 2.288294e-012, 1.850924e-012,
  0, 0, 0, 0,
  4.361411e-015, 3.241065e-015, 2.836004e-012, 4.089076e-012,
  0, 0, 0, 0,
  2.481924e-014, 4.588915e-015, 3.087062e-012, 3.97891e-012,
  0, 0, 0, 0,
  6.238681e-014, 1.317999e-014, 1.158023e-011, 1.6642e-011,
  0, 0, 0, 0,
  5.627758e-015, 9.417446e-015, 6.160226e-012, 1.108486e-011,
  0, 0, 0, 0,
  1.771642e-015, 2.680419e-015, 1.57823e-012, 2.112512e-012,
  0, 0, 0, 0,
  2.588279e-015, 4.118484e-015, 2.245029e-012, 3.227459e-012,
  0, 0, 0, 0,
  2.724948e-015, 3.016852e-015, 2.21635e-012, 2.116648e-012,
  0, 0, 0, 0,
  3.012183e-015, 2.661476e-015, 2.417814e-012, 3.473818e-012,
  0, 0, 0, 0,
  1.716797e-015, 2.104675e-015, 2.241525e-012, 2.08037e-012,
  0, 0, 0, 0,
  2.606593e-015, 2.413515e-015, 2.424249e-012, 2.662393e-012,
  0, 0, 0, 0,
  1.06685e-013, 1.849553e-014, 3.927916e-012, 5.386543e-012,
  0, 0, 0, 0,
  4.001445e-015, 4.976845e-015, 3.639199e-012, 4.827009e-012,
  0, 0, 0, 0,
  5.418235e-015, 1.764619e-014, 8.024574e-012, 1.672746e-011,
  0, 0, 0, 0,
  1.169177e-014, 2.254254e-014, 1.408532e-011, 2.710393e-011,
  0, 0, 0, 0,
  6.947993e-014, 1.364331e-014, 9.074936e-012, 1.723055e-011,
  0, 0, 0, 0,
  1.87749e-014, 4.442404e-015, 4.985761e-012, 7.179047e-012,
  0, 0, 0, 0,
  4.820141e-015, 3.764057e-015, 2.029939e-011, 2.096417e-011,
  0, 0, 0, 0,
  6.265568e-015, 3.18813e-015, 3.846894e-012, 5.783052e-012,
  0, 0, 0, 0,
  3.521326e-014, 6.088639e-015, 3.266785e-012, 4.475433e-012,
  0, 0, 0, 0,
  5.311318e-014, 8.571128e-015, 3.391036e-012, 3.746659e-012,
  0, 0, 0, 0,
  4.116185e-015, 3.247622e-015, 2.975418e-012, 3.87086e-012,
  0, 0, 0, 0,
  4.692993e-015, 2.49326e-015, 3.631151e-012, 4.5152e-012,
  0, 0, 0, 0,
  6.299499e-015, 7.161933e-015, 9.581882e-012, 1.603196e-011,
  0, 0, 0, 0,
  1.247087e-014, 2.816229e-014, 1.358628e-011, 2.447533e-011,
  0, 0, 0, 0,
  8.62653e-015, 2.621316e-014, 1.086534e-011, 2.024572e-011,
  0, 0, 0, 0,
  1.525159e-014, 2.064832e-014, 7.626642e-012, 1.665454e-011,
  0, 0, 0, 0,
  1.623171e-014, 1.614595e-014, 1.407585e-011, 1.867373e-011,
  0, 0, 0, 0,
  1.177632e-013, 2.73316e-014, 1.157627e-011, 1.993204e-011,
  0, 0, 0, 0,
  1.046535e-014, 1.359402e-014, 1.149396e-011, 1.757633e-011,
  0, 0, 0, 0,
  1.577483e-014, 1.421568e-014, 1.785454e-011, 2.599643e-011,
  0, 0, 0, 0,
  1.640491e-014, 2.548102e-014, 1.215365e-011, 2.565509e-011,
  0, 0, 0, 0,
  7.016225e-014, 2.466815e-014, 6.87008e-012, 1.131091e-011,
  0, 0, 0, 0,
  1.198414e-014, 1.888156e-014, 8.060902e-012, 1.487385e-011,
  0, 0, 0, 0,
  1.375827e-014, 1.507927e-014, 1.123364e-011, 2.113409e-011,
  0, 0, 0, 0,
  1.524937e-014, 2.523638e-014, 1.462058e-011, 1.984575e-011,
  0, 0, 0, 0,
  5.436518e-014, 2.926274e-014, 7.228724e-012, 1.516734e-011,
  0, 0, 0, 0,
  3.444709e-014, 3.475373e-014, 1.115428e-011, 2.517089e-011,
  0, 0, 0, 0,
  8.583998e-015, 1.616571e-014, 1.637789e-011, 2.226833e-011,
  0, 0, 0, 0,
  1.146147e-014, 8.790482e-015, 2.306914e-011, 2.577705e-011,
  0, 0, 0, 0,
  1.290497e-014, 1.418153e-014, 9.917366e-012, 1.930154e-011,
  0, 0, 0, 0,
  6.934389e-015, 2.27317e-014, 7.945472e-012, 1.553354e-011,
  0, 0, 0, 0,
  7.177606e-015, 4.325043e-015, 5.085519e-012, 7.049682e-012,
  0, 0, 0, 0,
  1.095103e-014, 9.001539e-015, 7.981267e-012, 1.254657e-011,
  0, 0, 0, 0,
  4.209247e-015, 1.78644e-014, 4.679371e-012, 1.213595e-011,
  0, 0, 0, 0,
  2.950632e-015, 7.493713e-015, 2.948726e-012, 4.624459e-012,
  0, 0, 0, 0,
  2.254945e-015, 3.82672e-015, 3.261793e-012, 3.619586e-012,
  0, 0, 0, 0,
  4.711707e-015, 1.981404e-014, 1.382152e-012, 2.161761e-012,
  0, 0, 0, 0,
  1.055566e-013, 2.089857e-014, 4.635874e-011, 7.250118e-011,
  0, 0, 0, 0,
  3.802581e-014, 1.09205e-014, 5.521834e-011, 7.028528e-011,
  0, 0, 0, 0,
  2.058163e-014, 3.018997e-014, 4.07851e-011, 3.693328e-011,
  0, 0, 0, 0,
  6.864524e-014, 7.283562e-014, 7.540268e-011, 1.158137e-010,
  0, 0, 0, 0,
  8.135063e-015, 6.60354e-015, 4.897068e-012, 5.754198e-012,
  0, 0, 0, 0,
  1.681889e-014, 2.531773e-014, 6.825181e-012, 1.292925e-011,
  0, 0, 0, 0,
  1.74432e-014, 2.341159e-014, 1.435865e-011, 2.909713e-011,
  0, 0, 0, 0,
  1.790694e-014, 3.393729e-014, 8.560984e-012, 2.114837e-011,
  0, 0, 0, 0,
  1.925109e-014, 1.186257e-014, 9.373782e-012, 1.928018e-011,
  0, 0, 0, 0,
  1.619991e-014, 1.061294e-014, 4.678054e-012, 8.118897e-012,
  0, 0, 0, 0,
  1.718749e-014, 1.182139e-014, 4.586677e-012, 7.961893e-012,
  0, 0, 0, 0,
  3.26894e-014, 9.238183e-015, 6.158051e-012, 1.054147e-011,
  0, 0, 0, 0,
  7.694454e-014, 1.835276e-014, 1.33191e-011, 2.78075e-011,
  0, 0, 0, 0,
  7.048926e-014, 1.571716e-014, 2.212943e-011, 3.213484e-011,
  0, 0, 0, 0,
  6.473966e-014, 1.645506e-014, 5.476353e-012, 1.253879e-011,
  0, 0, 0, 0,
  9.494933e-014, 3.918336e-014, 7.398771e-012, 2.166521e-011,
  0, 0, 0, 0,
  1.65369e-013, 4.321037e-014, 5.773822e-012, 2.3644e-011,
  0, 0, 0, 0,
  4.924805e-013, 8.698042e-014, 1.223866e-011, 5.27846e-011,
  0, 0, 0, 0,
  2.970196e-013, 6.499484e-014, 8.773607e-012, 3.099573e-011,
  0, 0, 0, 0,
  5.756564e-013, 1.134332e-013, 1.846443e-011, 6.036124e-011,
  0, 0, 0, 0,
  4.677106e-013, 1.249826e-013, 1.736266e-011, 6.039933e-011,
  0, 0, 0, 0,
  1.568357e-012, 3.166599e-013, 4.706868e-011, 2.120359e-010,
  0, 0, 0, 0,
  2.200924e-012, 4.542662e-013, 1.237609e-010, 4.473888e-010,
  0, 0, 0, 0,
  2.215381e-012, 4.5763e-013, 9.557223e-011, 3.543552e-010,
  0, 0, 0, 0,
  4.514672e-012, 1.231985e-012, 2.012716e-010, 8.07452e-010,
  0, 0, 0, 0,
  7.874095e-012, 2.308946e-012, 6.046839e-010, 1.780863e-009,
  0, 0, 0, 0,
  1.475921e-011, 4.483513e-012, 1.468548e-009, 7.386523e-009,
  0, 0, 0, 0,
  1.995111e-011, 5.154285e-012, 1.232016e-009, 4.745235e-009,
  0, 0, 0, 0,
  1.20035e-011, 4.192399e-012, 1.099677e-009, 3.569399e-009,
  0, 0, 0, 0,
  1.412768e-011, 4.25487e-012, 1.028984e-009, 3.526515e-009,
  0, 0, 0, 0,
  1.315001e-011, 4.849116e-012, 9.461839e-010, 3.716557e-009,
  0, 0, 0, 0,
  5.490014e-012, 2.269429e-012, 3.924493e-010, 1.594889e-009,
  0, 0, 0, 0,
  3.865434e-012, 9.624889e-013, 1.478686e-010, 6.4747e-010,
  0, 0, 0, 0,
  2.203305e-012, 5.872311e-013, 8.028886e-011, 3.250497e-010,
  0, 0, 0, 0,
  1.67064e-012, 4.465798e-013, 5.650126e-011, 2.423122e-010,
  0, 0, 0, 0,
  1.001771e-012, 2.212973e-013, 3.184522e-011, 1.355759e-010,
  0, 0, 0, 0,
  6.291355e-013, 2.060029e-013, 2.221619e-011, 7.471289e-011,
  0, 0, 0, 0,
  2.826256e-013, 1.904292e-013, 1.522798e-011, 6.10952e-011,
  0, 0, 0, 0,
  3.59502e-013, 2.108598e-013, 1.640569e-011, 6.440802e-011,
  0, 0, 0, 0,
  3.879068e-013, 8.418503e-014, 1.439835e-011, 4.311132e-011,
  0, 0, 0, 0,
  2.394185e-013, 6.473342e-014, 1.15589e-011, 1.978192e-011,
  0, 0, 0, 0,
  8.06509e-014, 4.422917e-014, 6.097193e-012, 1.618125e-011,
  0, 0, 0, 0,
  1.466545e-013, 4.29506e-014, 1.109481e-011, 2.449844e-011,
  0, 0, 0, 0,
  6.394536e-014, 2.99617e-014, 1.519262e-011, 3.350553e-011,
  0, 0, 0, 0,
  3.595593e-014, 2.912022e-014, 7.071106e-012, 1.855959e-011,
  0, 0, 0, 0,
  2.30986e-014, 2.740418e-014, 8.866859e-012, 1.638138e-011,
  0, 0, 0, 0,
  1.721929e-014, 3.864877e-014, 1.192653e-011, 2.519628e-011,
  0, 0, 0, 0,
  2.759351e-014, 3.349102e-014, 1.06533e-011, 2.623299e-011,
  0, 0, 0, 0,
  2.84056e-014, 1.927298e-014, 1.514664e-011, 2.746906e-011,
  0, 0, 0, 0,
  3.87148e-014, 3.421086e-014, 1.45773e-011, 2.798643e-011,
  0, 0, 0, 0,
  3.882149e-014, 6.555967e-014, 2.253514e-011, 3.341494e-011,
  0, 0, 0, 0,
  8.661633e-014, 4.289413e-014, 1.814356e-011, 4.177676e-011,
  0, 0, 0, 0,
  3.692772e-014, 4.389211e-014, 1.997741e-011, 3.004804e-011,
  0, 0, 0, 0,
  1.486962e-014, 2.725164e-014, 1.291623e-011, 2.56444e-011,
  0, 0, 0, 0,
  8.619712e-015, 3.266609e-014, 1.177327e-011, 2.642032e-011,
  0, 0, 0, 0,
  8.468478e-015, 2.205987e-014, 9.984764e-012, 1.917939e-011,
  0, 0, 0, 0,
  1.065547e-014, 2.892181e-014, 1.2091e-011, 2.596536e-011,
  0, 0, 0, 0,
  9.236548e-015, 2.624893e-014, 1.215079e-011, 1.949727e-011,
  0, 0, 0, 0,
  8.347152e-015, 3.342024e-014, 8.697055e-012, 1.847633e-011,
  0, 0, 0, 0,
  5.691599e-015, 2.685645e-014, 1.012772e-011, 2.309352e-011,
  0, 0, 0, 0,
  1.06684e-014, 2.18017e-014, 1.121389e-011, 2.280122e-011,
  0, 0, 0, 0,
  6.863783e-015, 3.482219e-014, 1.068965e-011, 2.233303e-011,
  0, 0, 0, 0,
  6.198883e-015, 2.987541e-014, 7.346093e-012, 1.715308e-011,
  0, 0, 0, 0,
  6.506812e-014, 4.624017e-014, 1.69319e-011, 3.415602e-011,
  0, 0, 0, 0,
  1.142922e-014, 5.286138e-014, 1.298065e-011, 2.390505e-011,
  0, 0, 0, 0,
  1.529704e-014, 3.191238e-014, 1.84358e-011, 3.033078e-011,
  0, 0, 0, 0,
  2.620135e-014, 3.078353e-014, 1.540137e-011, 2.72225e-011,
  0, 0, 0, 0,
  2.935503e-014, 8.915853e-014, 2.676522e-011, 6.877883e-011,
  0, 0, 0, 0,
  1.21707e-013, 5.585164e-014, 1.947591e-011, 3.580149e-011,
  0, 0, 0, 0,
  2.265289e-014, 5.293232e-014, 3.231048e-011, 6.396635e-011,
  0, 0, 0, 0,
  3.649415e-014, 5.206117e-014, 2.328022e-011, 5.145627e-011,
  0, 0, 0, 0,
  1.546747e-014, 4.022963e-014, 1.495096e-011, 3.300749e-011,
  0, 0, 0, 0,
  6.58983e-014, 3.676903e-014, 2.179031e-011, 4.625846e-011,
  0, 0, 0, 0,
  1.374733e-014, 2.551275e-014, 1.210293e-011, 2.472905e-011,
  0, 0, 0, 0,
  7.29188e-015, 3.327725e-014, 1.577065e-011, 3.457118e-011,
  0, 0, 0, 0,
  1.020532e-014, 3.77429e-014, 1.473799e-011, 2.67053e-011,
  0, 0, 0, 0,
  4.970964e-014, 3.038509e-014, 1.653028e-011, 2.702498e-011,
  0, 0, 0, 0,
  3.151747e-014, 4.452189e-014, 1.023111e-011, 1.963084e-011,
  0, 0, 0, 0,
  1.10471e-014, 3.365137e-014, 1.621116e-011, 3.256551e-011,
  0, 0, 0, 0,
  2.742757e-014, 2.770016e-014, 3.045984e-011, 3.890668e-011,
  0, 0, 0, 0,
  2.252682e-014, 3.518703e-014, 1.604133e-011, 3.174433e-011,
  0, 0, 0, 0,
  4.203568e-014, 6.020976e-014, 2.256444e-011, 4.241956e-011,
  0, 0, 0, 0,
  2.097828e-014, 9.851552e-014, 3.040372e-011, 5.860797e-011,
  0, 0, 0, 0,
  1.992231e-014, 3.508533e-014, 2.012633e-011, 3.989976e-011,
  0, 0, 0, 0,
  2.105902e-014, 7.100662e-014, 2.170214e-011, 4.194639e-011,
  0, 0, 0, 0,
  1.109858e-013, 5.175855e-014, 2.134019e-011, 3.818929e-011,
  0, 0, 0, 0,
  1.836377e-014, 4.957264e-014, 3.527409e-011, 6.371408e-011,
  0, 0, 0, 0,
  4.02174e-014, 5.912588e-014, 2.229784e-011, 4.83052e-011,
  0, 0, 0, 0,
  2.077174e-014, 6.506952e-014, 1.500026e-011, 4.02368e-011,
  0, 0, 0, 0,
  7.144949e-014, 2.918897e-014, 1.76122e-011, 4.218822e-011,
  0, 0, 0, 0,
  1.331252e-014, 3.189551e-014, 1.223883e-011, 2.066927e-011,
  0, 0, 0, 0,
  1.179943e-014, 2.457675e-014, 1.424397e-011, 3.387329e-011,
  0, 0, 0, 0,
  9.137475e-015, 3.030415e-014, 9.97327e-012, 2.018262e-011,
  0, 0, 0, 0,
  6.174616e-014, 3.213751e-014, 1.069398e-011, 2.25236e-011,
  0, 0, 0, 0,
  2.625371e-014, 3.464464e-014, 1.102186e-011, 2.553775e-011,
  0, 0, 0, 0,
  1.037509e-014, 2.679888e-014, 9.985872e-012, 2.258241e-011,
  0, 0, 0, 0,
  6.345648e-015, 2.877071e-014, 1.001488e-011, 1.978064e-011,
  0, 0, 0, 0,
  1.649697e-014, 2.685957e-014, 1.295954e-011, 3.146107e-011,
  0, 0, 0, 0,
  6.088275e-015, 1.908023e-014, 1.108876e-011, 2.098387e-011,
  0, 0, 0, 0,
  6.955451e-015, 1.488189e-014, 1.200924e-011, 2.735378e-011,
  0, 0, 0, 0,
  7.507749e-015, 3.037323e-014, 9.825082e-012, 1.960286e-011,
  0, 0, 0, 0,
  2.155788e-014, 6.004343e-014, 2.360921e-011, 4.039101e-011,
  0, 0, 0, 0,
  7.882885e-014, 4.277368e-014, 4.349025e-011, 7.001916e-011,
  0, 0, 0, 0,
  1.970126e-014, 5.134781e-014, 1.893855e-011, 3.30774e-011,
  0, 0, 0, 0,
  4.472265e-014, 9.474053e-014, 3.973658e-011, 6.76735e-011,
  0, 0, 0, 0,
  9.781154e-014, 8.039e-014, 4.745453e-011, 8.137306e-011,
  0, 0, 0, 0,
  9.013276e-014, 8.302256e-014, 2.864012e-011, 6.387533e-011,
  0, 0, 0, 0,
  7.672211e-014, 1.942086e-013, 5.45746e-011, 1.00564e-010,
  0, 0, 0, 0,
  1.136336e-013, 2.843811e-013, 1.698765e-010, 3.460537e-010,
  0, 0, 0, 0,
  1.070894e-013, 8.944199e-014, 7.379291e-011, 1.526747e-010,
  0, 0, 0, 0,
  1.512432e-013, 6.743794e-014, 8.429892e-011, 1.474175e-010,
  0, 0, 0, 0,
  9.320417e-014, 6.714283e-014, 6.673132e-011, 1.303355e-010,
  0, 0, 0, 0,
  2.345684e-013, 9.865169e-014, 1.894006e-010, 3.396697e-010,
  0, 0, 0, 0,
  1.885835e-013, 7.075345e-014, 1.587889e-010, 2.710367e-010,
  0, 0, 0, 0,
  1.762854e-013, 7.805764e-014, 1.803275e-010, 3.09266e-010,
  0, 0, 0, 0,
  1.513199e-013, 5.851996e-014, 1.178103e-010, 2.08872e-010,
  0, 0, 0, 0,
  3.143491e-013, 1.151426e-013, 2.906774e-010, 5.230142e-010,
  0, 0, 0, 0,
  7.726016e-014, 7.225127e-014, 8.383433e-011, 1.598848e-010,
  0, 0, 0, 0,
  1.348669e-013, 5.184281e-014, 8.509284e-011, 1.50553e-010,
  0, 0, 0, 0,
  8.041456e-014, 6.336793e-014, 3.410763e-011, 6.593719e-011,
  0, 0, 0, 0,
  7.139221e-014, 2.461746e-014, 3.022228e-011, 7.015959e-011,
  0, 0, 0, 0,
  4.745668e-014, 3.424171e-014, 3.187371e-011, 5.567076e-011,
  0, 0, 0, 0,
  2.777472e-014, 4.471226e-014, 2.75136e-011, 5.26203e-011,
  0, 0, 0, 0,
  1.093399e-013, 4.149273e-014, 4.376892e-011, 7.134332e-011,
  0, 0, 0, 0,
  4.699831e-014, 3.335677e-014, 2.885792e-011, 4.538788e-011,
  0, 0, 0, 0,
  2.567025e-014, 1.64673e-014, 1.42718e-011, 2.64362e-011,
  0, 0, 0, 0,
  2.107555e-014, 1.941502e-014, 1.415681e-011, 2.809876e-011,
  0, 0, 0, 0,
  3.072373e-014, 3.634558e-014, 2.111112e-011, 4.412745e-011,
  0, 0, 0, 0,
  2.997655e-014, 1.577344e-014, 1.369162e-011, 2.511175e-011,
  0, 0, 0, 0,
  2.041384e-014, 9.146818e-015, 8.434519e-012, 1.638784e-011,
  0, 0, 0, 0,
  9.371808e-015, 2.781115e-014, 1.128306e-011, 2.49562e-011,
  0, 0, 0, 0,
  5.419715e-014, 3.171895e-014, 1.321011e-011, 2.895399e-011,
  0, 0, 0, 0,
  3.547946e-014, 3.672922e-014, 2.154337e-011, 4.925265e-011,
  0, 0, 0, 0,
  2.593198e-014, 5.039267e-014, 1.970452e-011, 3.92941e-011,
  0, 0, 0, 0,
  2.476785e-014, 4.100809e-014, 2.11725e-011, 3.234048e-011,
  0, 0, 0, 0,
  3.392948e-014, 1.874824e-014, 2.13699e-011, 3.641557e-011,
  0, 0, 0, 0,
  7.17803e-014, 3.724518e-014, 2.895099e-011, 5.691797e-011,
  0, 0, 0, 0,
  1.160269e-013, 6.473234e-014, 6.678892e-011, 1.165414e-010,
  0, 0, 0, 0,
  7.717155e-014, 3.534261e-014, 5.679513e-011, 1.023546e-010,
  0, 0, 0, 0,
  6.293869e-014, 4.554737e-014, 3.784369e-011, 6.880013e-011,
  0, 0, 0, 0,
  5.05885e-014, 4.580615e-014, 4.681253e-011, 6.858519e-011,
  0, 0, 0, 0,
  7.709478e-014, 2.909885e-014, 6.217439e-011, 1.081382e-010,
  0, 0, 0, 0,
  4.405264e-014, 2.091635e-014, 3.767049e-011, 7.628538e-011,
  0, 0, 0, 0,
  9.018699e-014, 3.880102e-014, 8.598853e-011, 1.549407e-010,
  0, 0, 0, 0,
  1.364967e-013, 4.546036e-014, 1.097722e-010, 2.149158e-010,
  0, 0, 0, 0,
  8.828309e-014, 5.230945e-014, 8.373791e-011, 1.601883e-010,
  0, 0, 0, 0,
  1.302017e-013, 5.375077e-014, 1.279537e-010, 2.387478e-010,
  0, 0, 0, 0,
  1.359995e-013, 5.994391e-014, 1.493419e-010, 2.715138e-010,
  0, 0, 0, 0,
  6.028554e-013, 1.263288e-013, 8.11229e-010, 1.470276e-009,
  0, 0, 0, 0,
  1.125597e-013, 1.055422e-013, 1.178942e-010, 2.173885e-010,
  0, 0, 0, 0,
  1.045356e-013, 5.347118e-014, 1.234026e-010, 2.18707e-010,
  0, 0, 0, 0,
  1.57017e-013, 6.123134e-014, 1.902516e-010, 3.589443e-010,
  0, 0, 0, 0,
  3.395826e-013, 9.514426e-014, 3.916099e-010, 7.186109e-010,
  0, 0, 0, 0,
  1.464212e-013, 4.096306e-014, 1.37371e-010, 2.577979e-010,
  0, 0, 0, 0,
  1.424627e-013, 5.231555e-014, 1.22805e-010, 2.308277e-010,
  0, 0, 0, 0,
  6.341962e-014, 5.002268e-014, 4.175249e-011, 7.289843e-011,
  0, 0, 0, 0,
  7.771924e-014, 4.917626e-014, 8.071489e-011, 1.506262e-010,
  0, 0, 0, 0,
  1.000808e-013, 3.726718e-014, 2.296875e-011, 3.990439e-011,
  0, 0, 0, 0,
  4.28843e-014, 5.631919e-014, 3.336018e-011, 6.838542e-011,
  0, 0, 0, 0,
  4.047212e-014, 2.440971e-014, 2.261095e-011, 4.71806e-011,
  0, 0, 0, 0,
  6.044769e-014, 3.477121e-014, 2.57975e-011, 5.036619e-011,
  0, 0, 0, 0,
  8.991615e-014, 4.531227e-014, 2.188898e-011, 4.451266e-011,
  0, 0, 0, 0,
  3.634398e-014, 2.778426e-014, 2.762787e-011, 5.473272e-011,
  0, 0, 0, 0,
  6.672326e-014, 4.025913e-014, 3.491484e-011, 6.704241e-011,
  0, 0, 0, 0,
  1.775226e-013, 1.317629e-013, 1.034723e-010, 1.947185e-010,
  0, 0, 0, 0,
  9.870152e-014, 4.226493e-014, 8.984304e-011, 1.707961e-010,
  0, 0, 0, 0,
  5.440962e-014, 6.154058e-014, 4.743817e-011, 8.754662e-011,
  0, 0, 0, 0,
  6.565524e-014, 8.784221e-014, 4.157865e-011, 7.827487e-011,
  0, 0, 0, 0,
  1.165728e-013, 9.545077e-014, 7.418069e-011, 1.45987e-010,
  0, 0, 0, 0,
  9.529317e-014, 6.57568e-014, 1.018813e-010, 1.900145e-010,
  0, 0, 0, 0,
  1.002961e-013, 6.526004e-014, 6.456384e-011, 1.183931e-010,
  0, 0, 0, 0,
  8.028459e-014, 4.582333e-014, 5.649537e-011, 9.071962e-011,
  0, 0, 0, 0,
  7.342647e-014, 5.130386e-014, 5.011123e-011, 9.465406e-011,
  0, 0, 0, 0,
  7.857214e-014, 4.58865e-014, 6.283212e-011, 9.773007e-011,
  0, 0, 0, 0,
  8.83905e-014, 5.414277e-014, 3.467389e-011, 6.828177e-011,
  0, 0, 0, 0,
  7.444716e-014, 4.266048e-014, 4.564492e-011, 8.227702e-011,
  0, 0, 0, 0,
  9.047282e-014, 6.316378e-014, 5.567314e-011, 9.909344e-011,
  0, 0, 0, 0,
  9.264485e-014, 4.883122e-014, 6.050219e-011, 1.021559e-010,
  0, 0, 0, 0,
  9.850919e-014, 4.139415e-014, 3.836365e-011, 6.638814e-011,
  0, 0, 0, 0,
  3.599612e-014, 3.240765e-014, 3.491587e-011, 6.70835e-011,
  0, 0, 0, 0,
  3.754406e-014, 2.969865e-014, 2.635723e-011, 4.94439e-011,
  0, 0, 0, 0,
  3.640988e-014, 2.868619e-014, 2.824295e-011, 4.943968e-011,
  0, 0, 0, 0,
  5.230357e-014, 4.49596e-014, 3.786865e-011, 7.585792e-011,
  0, 0, 0, 0,
  7.833351e-014, 4.122366e-014, 4.519893e-011, 8.313344e-011,
  0, 0, 0, 0,
  5.039737e-014, 4.214708e-014, 3.984737e-011, 6.613955e-011,
  0, 0, 0, 0,
  8.168549e-014, 5.128204e-014, 7.11271e-011, 1.265354e-010,
  0, 0, 0, 0,
  1.068711e-013, 4.913208e-014, 5.943027e-011, 1.13152e-010,
  0, 0, 0, 0,
  1.205275e-013, 5.094323e-014, 1.094955e-010, 2.008561e-010,
  0, 0, 0, 0,
  2.668903e-013, 9.350824e-014, 2.413332e-010, 4.52833e-010,
  0, 0, 0, 0,
  3.544602e-013, 9.652883e-014, 4.591514e-010, 8.786151e-010,
  0, 0, 0, 0,
  1.858288e-013, 4.405114e-014, 2.203927e-010, 3.97249e-010,
  0, 0, 0, 0,
  2.388443e-013, 7.86612e-014, 2.542462e-010, 4.724706e-010,
  0, 0, 0, 0,
  3.63674e-013, 8.662284e-014, 4.384403e-010, 8.240879e-010,
  0, 0, 0, 0,
  1.935988e-013, 7.943513e-014, 1.877663e-010, 3.527481e-010,
  0, 0, 0, 0,
  3.145616e-013, 9.679144e-014, 2.637674e-010, 5.032745e-010,
  0, 0, 0, 0,
  7.352571e-014, 3.29291e-014, 6.827021e-011, 1.149723e-010,
  0, 0, 0, 0,
  9.986404e-014, 4.921821e-014, 8.804293e-011, 1.461863e-010,
  0, 0, 0, 0,
  7.28696e-014, 4.379705e-014, 4.257348e-011, 6.963503e-011,
  0, 0, 0, 0,
  1.625041e-013, 8.015596e-014, 1.697229e-010, 3.03277e-010,
  0, 0, 0, 0,
  8.361589e-014, 5.978884e-014, 6.605736e-011, 1.232189e-010,
  0, 0, 0, 0,
  7.73223e-014, 3.79942e-014, 6.786013e-011, 1.166166e-010,
  0, 0, 0, 0,
  9.547993e-014, 5.627743e-014, 6.029409e-011, 1.218185e-010,
  0, 0, 0, 0,
  8.833099e-014, 3.439404e-014, 5.651541e-011, 9.961838e-011,
  0, 0, 0, 0,
  1.395841e-013, 5.164294e-014, 9.279456e-011, 1.558533e-010,
  0, 0, 0, 0,
  8.621526e-014, 4.201749e-014, 6.081853e-011, 1.239718e-010,
  0, 0, 0, 0,
  1.203116e-013, 5.557703e-014, 7.746309e-011, 1.346355e-010,
  0, 0, 0, 0,
  1.462693e-013, 5.19615e-014, 7.585181e-011, 1.367135e-010,
  0, 0, 0, 0,
  1.164377e-013, 6.167779e-014, 6.776116e-011, 1.268826e-010,
  0, 0, 0, 0,
  1.54322e-013, 7.066996e-014, 1.14183e-010, 2.137713e-010,
  0, 0, 0, 0,
  1.892204e-013, 7.881664e-014, 1.731257e-010, 3.161582e-010,
  0, 0, 0, 0,
  1.98654e-013, 1.237774e-013, 2.109916e-010, 3.864092e-010,
  0, 0, 0, 0,
  1.584657e-013, 9.736016e-014, 2.024889e-010, 3.888563e-010,
  0, 0, 0, 0,
  3.026807e-013, 1.172425e-013, 3.885393e-010, 7.379104e-010,
  0, 0, 0, 0,
  2.921683e-013, 1.022868e-013, 3.813279e-010, 7.168287e-010,
  0, 0, 0, 0,
  4.210753e-013, 1.116401e-013, 6.140866e-010, 1.119784e-009,
  0, 0, 0, 0,
  3.634091e-013, 1.074401e-013, 4.452703e-010, 8.126159e-010,
  0, 0, 0, 0,
  8.245219e-015, 2.749391e-015, 5.924504e-012, 8.914372e-012,
  0, 0, 0, 0,
  2.821222e-014, 5.1217e-015, 3.308528e-011, 2.845982e-011,
  0, 0, 0, 0,
  9.389708e-014, 1.502664e-014, 7.393883e-012, 7.437385e-012,
  0, 0, 0, 0,
  7.40097e-015, 1.447214e-014, 8.055376e-012, 8.503475e-012,
  0, 0, 0, 0,
  5.701586e-015, 8.577961e-015, 4.898344e-012, 5.498971e-012,
  0, 0, 0, 0,
  6.664415e-015, 4.738753e-015, 1.238156e-011, 2.094718e-011,
  0, 0, 0, 0,
  8.236792e-014, 1.436028e-014, 9.706983e-012, 1.350546e-011,
  0, 0, 0, 0,
  4.758336e-015, 1.96338e-014, 9.173566e-012, 1.812147e-011,
  0, 0, 0, 0,
  3.497361e-014, 8.412591e-015, 3.701432e-011, 4.443189e-011,
  0, 0, 0, 0,
  4.150787e-014, 1.80558e-013, 3.456206e-011, 4.282961e-011,
  0, 0, 0, 0,
  8.279759e-014, 1.567113e-014, 8.374341e-012, 1.080986e-011,
  0, 0, 0, 0,
  9.881461e-015, 4.270716e-015, 3.409273e-012, 4.682282e-012,
  0, 0, 0, 0,
  4.76025e-015, 4.081437e-015, 8.945727e-012, 9.454428e-012,
  0, 0, 0, 0,
  1.217823e-014, 2.967355e-015, 8.984484e-012, 1.209882e-011,
  0, 0, 0, 0,
  8.153581e-015, 2.415399e-015, 4.10582e-012, 6.639279e-012,
  0, 0, 0, 0,
  9.854083e-015, 3.059465e-015, 9.382503e-012, 1.537318e-011,
  0, 0, 0, 0,
  3.831667e-014, 7.521022e-015, 2.736477e-011, 4.798282e-011,
  0, 0, 0, 0,
  4.937596e-015, 2.174168e-015, 4.919064e-012, 7.84401e-012,
  0, 0, 0, 0,
  6.231729e-015, 1.094212e-014, 4.937712e-012, 8.095478e-012,
  0, 0, 0, 0,
  9.628898e-015, 7.164772e-015, 9.027606e-012, 1.53515e-011,
  0, 0, 0, 0,
  1.372369e-014, 3.354389e-015, 1.152143e-011, 1.820731e-011,
  0, 0, 0, 0,
  8.548906e-015, 2.991607e-015, 6.226562e-012, 8.934128e-012,
  0, 0, 0, 0,
  3.693211e-014, 6.711114e-015, 2.195857e-011, 3.848161e-011,
  0, 0, 0, 0,
  9.777824e-014, 1.597997e-014, 2.19448e-011, 3.57174e-011,
  0, 0, 0, 0,
  1.121175e-014, 6.712264e-015, 7.392597e-012, 1.126128e-011,
  0, 0, 0, 0,
  4.604358e-015, 4.407306e-015, 7.579196e-012, 9.224741e-012,
  0, 0, 0, 0,
  1.741945e-014, 7.317899e-015, 1.002804e-011, 1.91927e-011,
  0, 0, 0, 0,
  9.449142e-014, 1.490171e-014, 2.182265e-011, 2.85392e-011,
  0, 0, 0, 0,
  9.980078e-015, 4.684251e-015, 6.705341e-012, 1.107942e-011,
  0, 0, 0, 0,
  9.531693e-015, 3.331888e-015, 8.668294e-012, 1.397604e-011,
  0, 0, 0, 0,
  3.532102e-015, 2.617257e-015, 3.300042e-012, 2.965596e-012,
  0, 0, 0, 0,
  1.043838e-014, 4.421468e-015, 8.392126e-012, 2.142988e-011,
  0, 0, 0, 0,
  1.352404e-014, 3.142751e-015, 1.047925e-011, 1.851302e-011,
  0, 0, 0, 0,
  1.506098e-014, 3.172121e-015, 4.826817e-012, 1.090604e-011,
  0, 0, 0, 0,
  7.796133e-015, 3.705328e-015, 8.593553e-012, 1.009749e-011,
  0, 0, 0, 0,
  6.328239e-014, 1.067984e-014, 5.950705e-012, 7.830203e-012,
  0, 0, 0, 0,
  7.463913e-014, 1.209211e-014, 2.776504e-011, 4.543091e-011,
  0, 0, 0, 0,
  1.184054e-014, 3.035333e-015, 5.107253e-012, 7.954153e-012,
  0, 0, 0, 0,
  7.141414e-015, 2.714262e-015, 3.213292e-012, 4.022485e-012,
  0, 0, 0, 0,
  1.416925e-014, 3.474648e-015, 2.086592e-012, 3.144362e-012,
  0, 0, 0, 0,
  7.214404e-014, 1.176398e-014, 2.366699e-012, 4.278234e-012,
  0, 0, 0, 0,
  2.806959e-014, 5.41719e-015, 1.122988e-011, 2.078683e-011,
  0, 0, 0, 0,
  8.935019e-015, 3.901524e-015, 4.958502e-012, 8.202606e-012,
  0, 0, 0, 0,
  5.079515e-015, 3.76619e-015, 3.477586e-012, 6.318739e-012,
  0, 0, 0, 0,
  9.052874e-014, 1.422931e-014, 3.003449e-012, 3.943445e-012,
  0, 0, 0, 0,
  6.285231e-015, 4.776241e-015, 3.300233e-012, 3.952255e-012,
  0, 0, 0, 0,
  4.955287e-015, 1.721816e-014, 4.012582e-012, 1.06097e-011,
  0, 0, 0, 0,
  4.91665e-015, 8.585477e-015, 3.90548e-012, 6.131949e-012,
  0, 0, 0, 0,
  1.18645e-013, 3.334048e-014, 1.132488e-011, 2.123727e-011,
  0, 0, 0, 0,
  1.914977e-014, 5.017095e-015, 2.266067e-011, 2.607829e-011,
  0, 0, 0, 0,
  4.834108e-015, 3.201082e-015, 2.525033e-012, 2.890519e-012,
  0, 0, 0, 0,
  2.563232e-015, 2.047505e-015, 2.524198e-012, 2.011981e-012,
  0, 0, 0, 0,
  4.56681e-014, 7.968329e-015, 2.774859e-012, 4.292083e-012,
  0, 0, 0, 0,
  3.577797e-014, 6.635783e-015, 4.377601e-012, 6.184519e-012,
  0, 0, 0, 0,
  3.221164e-015, 2.253525e-015, 2.91521e-012, 3.293924e-012,
  0, 0, 0, 0,
  5.527321e-015, 2.853318e-015, 2.935014e-012, 4.513733e-012,
  0, 0, 0, 0,
  2.531723e-014, 5.231446e-015, 6.730198e-012, 8.831937e-012,
  0, 0, 0, 0,
  6.317815e-014, 1.18416e-014, 1.263384e-011, 1.996874e-011,
  0, 0, 0, 0,
  4.650762e-015, 6.829332e-015, 4.774773e-012, 7.807204e-012,
  0, 0, 0, 0,
  3.005481e-015, 2.617012e-015, 1.985854e-012, 2.330675e-012,
  0, 0, 0, 0,
  2.942687e-015, 2.047573e-015, 2.658781e-012, 2.403037e-012,
  0, 0, 0, 0,
  2.480497e-015, 2.364422e-015, 1.613827e-012, 1.580827e-012,
  0, 0, 0, 0,
  3.031845e-015, 2.616277e-015, 2.743387e-012, 3.640604e-012,
  0, 0, 0, 0,
  3.038936e-015, 3.171663e-015, 1.542971e-012, 2.251698e-012,
  0, 0, 0, 0,
  2.262437e-015, 2.257719e-015, 1.548836e-012, 1.407619e-012,
  0, 0, 0, 0,
  1.188441e-013, 2.3497e-014, 2.310627e-012, 4.369702e-012,
  0, 0, 0, 0,
  4.646952e-015, 5.574886e-015, 1.978826e-012, 2.935514e-012,
  0, 0, 0, 0,
  3.654404e-015, 1.290466e-014, 5.243851e-012, 8.904322e-012,
  0, 0, 0, 0,
  6.596664e-015, 1.319522e-014, 7.518763e-012, 1.205019e-011,
  0, 0, 0, 0,
  6.937083e-014, 1.133716e-014, 5.757798e-012, 1.14841e-011,
  0, 0, 0, 0,
  1.969442e-014, 3.823595e-015, 3.613679e-012, 5.246633e-012,
  0, 0, 0, 0,
  3.993058e-015, 4.731704e-015, 2.151803e-011, 2.292826e-011,
  0, 0, 0, 0,
  6.984075e-015, 2.584689e-015, 6.141975e-012, 1.012516e-011,
  0, 0, 0, 0,
  3.640612e-014, 6.382724e-015, 3.390796e-012, 3.977046e-012,
  0, 0, 0, 0,
  5.298883e-014, 8.463912e-015, 4.379013e-012, 7.752683e-012,
  0, 0, 0, 0,
  4.51099e-015, 2.669397e-015, 3.613032e-012, 6.017157e-012,
  0, 0, 0, 0,
  7.126524e-015, 3.749868e-015, 4.578807e-012, 6.137025e-012,
  0, 0, 0, 0,
  1.610687e-014, 5.717206e-015, 1.52756e-011, 2.37563e-011,
  0, 0, 0, 0,
  2.699114e-014, 1.120592e-014, 2.598642e-011, 4.126147e-011,
  0, 0, 0, 0,
  1.000906e-014, 1.083093e-014, 6.96212e-012, 1.296023e-011,
  0, 0, 0, 0,
  1.364959e-014, 7.93018e-015, 1.237451e-011, 2.12724e-011,
  0, 0, 0, 0,
  2.305524e-014, 1.273999e-014, 1.604136e-011, 3.21585e-011,
  0, 0, 0, 0,
  1.228574e-013, 2.195423e-014, 9.776244e-012, 1.089954e-011,
  0, 0, 0, 0,
  2.887105e-014, 1.194441e-014, 2.300502e-011, 4.341406e-011,
  0, 0, 0, 0,
  1.964813e-014, 1.139767e-014, 1.620887e-011, 2.778422e-011,
  0, 0, 0, 0,
  1.331339e-014, 1.407523e-014, 1.492811e-011, 2.217625e-011,
  0, 0, 0, 0,
  7.606449e-014, 1.600668e-014, 8.349162e-012, 1.271726e-011,
  0, 0, 0, 0,
  1.288618e-014, 1.164023e-014, 7.721922e-012, 1.25672e-011,
  0, 0, 0, 0,
  1.572167e-014, 1.505653e-014, 1.035208e-011, 1.704535e-011,
  0, 0, 0, 0,
  1.8295e-014, 3.571938e-014, 1.638269e-011, 1.918662e-011,
  0, 0, 0, 0,
  5.335799e-014, 2.226933e-014, 8.659787e-012, 1.106163e-011,
  0, 0, 0, 0,
  3.379098e-014, 1.475951e-014, 6.886161e-012, 9.672007e-012,
  0, 0, 0, 0,
  1.566645e-014, 2.079346e-014, 1.143797e-011, 2.338241e-011,
  0, 0, 0, 0,
  1.590012e-014, 8.029393e-015, 2.209324e-011, 2.49223e-011,
  0, 0, 0, 0,
  2.068637e-014, 1.288773e-014, 8.445875e-012, 1.959003e-011,
  0, 0, 0, 0,
  5.832519e-015, 1.339964e-014, 7.264235e-012, 1.029658e-011,
  0, 0, 0, 0,
  9.08535e-015, 3.519063e-015, 7.428358e-012, 1.31577e-011,
  0, 0, 0, 0,
  1.024318e-014, 6.490899e-015, 6.413928e-012, 1.050671e-011,
  0, 0, 0, 0,
  5.511369e-015, 4.389578e-015, 4.050405e-012, 8.915253e-012,
  0, 0, 0, 0,
  4.857765e-015, 3.217433e-015, 2.788038e-012, 2.873782e-012,
  0, 0, 0, 0,
  3.48909e-015, 4.206863e-015, 2.219022e-012, 2.036361e-012,
  0, 0, 0, 0,
  6.149559e-015, 2.056386e-014, 2.498811e-012, 2.165892e-012,
  0, 0, 0, 0,
  1.204007e-013, 2.033228e-014, 4.805512e-011, 8.859792e-011,
  0, 0, 0, 0,
  9.355064e-014, 1.707255e-014, 8.880002e-011, 1.247027e-010,
  0, 0, 0, 0,
  5.149099e-014, 1.389959e-014, 4.830325e-011, 6.184914e-011,
  0, 0, 0, 0,
  2.259922e-013, 4.701381e-014, 1.302523e-010, 2.128456e-010,
  0, 0, 0, 0,
  5.317712e-015, 6.065603e-015, 3.983781e-012, 7.180753e-012,
  0, 0, 0, 0,
  1.479351e-014, 9.438992e-015, 7.889967e-012, 1.68282e-011,
  0, 0, 0, 0,
  6.618882e-014, 2.433619e-014, 5.768174e-011, 1.061984e-010,
  0, 0, 0, 0,
  1.664855e-014, 1.367018e-014, 5.454358e-012, 1.314981e-011,
  0, 0, 0, 0,
  1.221156e-014, 9.842314e-015, 1.13018e-011, 1.970288e-011,
  0, 0, 0, 0,
  1.071614e-014, 4.363382e-015, 4.178729e-012, 4.843178e-012,
  0, 0, 0, 0,
  1.811851e-014, 6.838268e-015, 3.765973e-012, 8.470701e-012,
  0, 0, 0, 0,
  3.213205e-014, 7.018306e-015, 3.317712e-012, 9.84011e-012,
  0, 0, 0, 0,
  7.477559e-014, 1.380472e-014, 1.400058e-011, 3.458109e-011,
  0, 0, 0, 0,
  6.042774e-014, 1.444956e-014, 3.424157e-011, 4.432908e-011,
  0, 0, 0, 0,
  4.427815e-014, 1.309407e-014, 3.793661e-012, 1.211115e-011,
  0, 0, 0, 0,
  6.144027e-014, 1.723548e-014, 6.355529e-012, 1.464055e-011,
  0, 0, 0, 0,
  1.628697e-013, 4.339134e-014, 5.978134e-012, 2.541528e-011,
  0, 0, 0, 0,
  3.995689e-013, 7.127904e-014, 9.015504e-012, 4.842295e-011,
  0, 0, 0, 0,
  2.936346e-013, 6.421864e-014, 8.617512e-012, 3.777573e-011,
  0, 0, 0, 0,
  6.026803e-013, 1.106405e-013, 1.777827e-011, 8.725165e-011,
  0, 0, 0, 0,
  6.788173e-013, 1.37456e-013, 1.846509e-011, 7.986727e-011,
  0, 0, 0, 0,
  1.658069e-012, 3.287325e-013, 5.242927e-011, 2.239006e-010,
  0, 0, 0, 0,
  2.467965e-012, 4.995194e-013, 1.378083e-010, 4.979411e-010,
  0, 0, 0, 0,
  2.337737e-012, 5.626699e-013, 1.036892e-010, 3.964575e-010,
  0, 0, 0, 0,
  3.961989e-012, 1.191232e-012, 1.861697e-010, 7.264769e-010,
  0, 0, 0, 0,
  9.349069e-012, 2.505017e-012, 7.11377e-010, 1.92214e-009,
  0, 0, 0, 0,
  1.481136e-011, 4.511911e-012, 1.443473e-009, 7.259866e-009,
  0, 0, 0, 0,
  2.032163e-011, 5.676453e-012, 1.298993e-009, 4.581221e-009,
  0, 0, 0, 0,
  1.355657e-011, 4.322091e-012, 1.096166e-009, 3.749166e-009,
  0, 0, 0, 0,
  1.646265e-011, 5.264011e-012, 1.22713e-009, 4.123655e-009,
  0, 0, 0, 0,
  1.382944e-011, 5.73432e-012, 1.200781e-009, 4.779837e-009,
  0, 0, 0, 0,
  4.901115e-012, 2.223143e-012, 3.892829e-010, 1.578622e-009,
  0, 0, 0, 0,
  3.989835e-012, 8.83118e-013, 1.551417e-010, 6.87405e-010,
  0, 0, 0, 0,
  2.138249e-012, 5.257985e-013, 7.452472e-011, 3.216811e-010,
  0, 0, 0, 0,
  1.978716e-012, 5.719653e-013, 5.994173e-011, 2.93346e-010,
  0, 0, 0, 0,
  1.151161e-012, 3.761426e-013, 4.737695e-011, 1.626222e-010,
  0, 0, 0, 0,
  5.519713e-013, 2.882669e-013, 2.203374e-011, 7.773058e-011,
  0, 0, 0, 0,
  3.638843e-013, 2.79434e-013, 1.915435e-011, 5.465074e-011,
  0, 0, 0, 0,
  4.11433e-013, 2.492498e-013, 1.721525e-011, 5.373434e-011,
  0, 0, 0, 0,
  2.421465e-013, 7.879702e-014, 1.5236e-011, 4.815837e-011,
  0, 0, 0, 0,
  2.913844e-013, 6.242787e-014, 9.544946e-012, 2.777384e-011,
  0, 0, 0, 0,
  8.326967e-014, 2.859127e-014, 6.914312e-012, 1.881826e-011,
  0, 0, 0, 0,
  1.143928e-013, 3.029438e-014, 8.993173e-012, 2.965332e-011,
  0, 0, 0, 0,
  6.151831e-014, 8.118372e-014, 2.019253e-011, 4.31822e-011,
  0, 0, 0, 0,
  3.217766e-014, 2.613587e-014, 8.733306e-012, 1.57972e-011,
  0, 0, 0, 0,
  2.517223e-014, 3.171766e-014, 1.515754e-011, 4.259883e-011,
  0, 0, 0, 0,
  2.468978e-014, 2.769486e-014, 1.318049e-011, 3.244897e-011,
  0, 0, 0, 0,
  2.667213e-014, 4.692548e-014, 1.518481e-011, 2.305488e-011,
  0, 0, 0, 0,
  3.602592e-014, 3.634007e-014, 2.038219e-011, 4.488279e-011,
  0, 0, 0, 0,
  1.012867e-013, 6.3016e-014, 3.610001e-011, 6.785175e-011,
  0, 0, 0, 0,
  4.254195e-014, 6.032405e-014, 2.532274e-011, 6.878701e-011,
  0, 0, 0, 0,
  8.355174e-014, 5.695599e-014, 1.740548e-011, 3.349981e-011,
  0, 0, 0, 0,
  2.868618e-014, 5.624633e-014, 2.686656e-011, 5.344817e-011,
  0, 0, 0, 0,
  3.481717e-014, 3.77053e-014, 2.128956e-011, 4.887673e-011,
  0, 0, 0, 0,
  1.219019e-014, 3.48972e-014, 1.156091e-011, 2.710094e-011,
  0, 0, 0, 0,
  9.955659e-015, 3.057048e-014, 1.621393e-011, 3.918798e-011,
  0, 0, 0, 0,
  9.246334e-015, 3.301143e-014, 1.083911e-011, 2.830699e-011,
  0, 0, 0, 0,
  9.597608e-015, 2.524576e-014, 1.645918e-011, 1.695272e-011,
  0, 0, 0, 0,
  6.671157e-015, 1.320952e-014, 6.724732e-012, 1.619649e-011,
  0, 0, 0, 0,
  7.162367e-015, 3.336572e-014, 1.047294e-011, 1.887736e-011,
  0, 0, 0, 0,
  6.48096e-015, 1.767205e-014, 6.5704e-012, 1.373e-011,
  0, 0, 0, 0,
  7.802856e-015, 3.165209e-014, 8.610284e-012, 1.58382e-011,
  0, 0, 0, 0,
  6.296983e-015, 3.155348e-014, 8.16633e-012, 1.56001e-011,
  0, 0, 0, 0,
  2.996286e-014, 5.15985e-014, 2.807257e-011, 5.462844e-011,
  0, 0, 0, 0,
  9.556824e-015, 5.054889e-014, 1.43799e-011, 3.108588e-011,
  0, 0, 0, 0,
  1.326974e-014, 3.257912e-014, 1.295119e-011, 2.533073e-011,
  0, 0, 0, 0,
  2.982429e-014, 6.712358e-014, 3.72618e-011, 7.649387e-011,
  0, 0, 0, 0,
  2.445026e-014, 8.513661e-014, 3.473799e-011, 6.88532e-011,
  0, 0, 0, 0,
  1.232498e-013, 6.08487e-014, 2.987844e-011, 5.43402e-011,
  0, 0, 0, 0,
  2.260036e-014, 7.869633e-014, 4.034547e-011, 7.696978e-011,
  0, 0, 0, 0,
  3.032457e-014, 6.024482e-014, 2.931784e-011, 5.740292e-011,
  0, 0, 0, 0,
  1.626784e-014, 6.593392e-014, 2.052262e-011, 4.189971e-011,
  0, 0, 0, 0,
  6.789493e-014, 5.01945e-014, 1.305046e-011, 3.829973e-011,
  0, 0, 0, 0,
  1.519971e-014, 3.031838e-014, 1.76025e-011, 4.146792e-011,
  0, 0, 0, 0,
  8.477526e-015, 4.0457e-014, 1.291299e-011, 3.309748e-011,
  0, 0, 0, 0,
  1.297802e-014, 4.808899e-014, 1.918245e-011, 3.612212e-011,
  0, 0, 0, 0,
  4.888648e-014, 5.63435e-014, 1.677989e-011, 4.449636e-011,
  0, 0, 0, 0,
  3.40104e-014, 6.611757e-014, 1.302208e-011, 3.019807e-011,
  0, 0, 0, 0,
  1.360018e-014, 5.845023e-014, 1.412393e-011, 3.120622e-011,
  0, 0, 0, 0,
  2.720743e-014, 5.026153e-014, 3.852611e-011, 7.270477e-011,
  0, 0, 0, 0,
  2.39267e-014, 6.877956e-014, 1.618373e-011, 3.926049e-011,
  0, 0, 0, 0,
  2.44986e-014, 5.468774e-014, 2.550606e-011, 5.213269e-011,
  0, 0, 0, 0,
  2.643949e-014, 4.995571e-014, 3.269434e-011, 7.555329e-011,
  0, 0, 0, 0,
  2.433027e-014, 7.104648e-014, 1.572444e-011, 3.20798e-011,
  0, 0, 0, 0,
  2.243127e-014, 7.158447e-014, 2.259992e-011, 3.930001e-011,
  0, 0, 0, 0,
  1.241049e-013, 6.523148e-014, 2.968926e-011, 5.782112e-011,
  0, 0, 0, 0,
  3.728947e-014, 9.10857e-014, 3.508129e-011, 7.436375e-011,
  0, 0, 0, 0,
  3.524473e-014, 8.75486e-014, 3.103234e-011, 7.707314e-011,
  0, 0, 0, 0,
  1.3712e-014, 6.235067e-014, 2.109861e-011, 5.084574e-011,
  0, 0, 0, 0,
  7.338845e-014, 4.940115e-014, 9.976671e-012, 2.616044e-011,
  0, 0, 0, 0,
  1.770045e-014, 3.725108e-014, 1.839296e-011, 4.120796e-011,
  0, 0, 0, 0,
  1.817725e-014, 4.561646e-014, 1.803432e-011, 3.823186e-011,
  0, 0, 0, 0,
  1.27037e-014, 3.261563e-014, 1.615763e-011, 4.186289e-011,
  0, 0, 0, 0,
  6.308481e-014, 2.807762e-014, 7.955081e-012, 1.949222e-011,
  0, 0, 0, 0,
  2.215606e-014, 1.876635e-014, 9.412641e-012, 1.79901e-011,
  0, 0, 0, 0,
  1.148692e-014, 2.366245e-014, 1.071953e-011, 2.427576e-011,
  0, 0, 0, 0,
  7.378244e-015, 2.179012e-014, 8.299229e-012, 1.931561e-011,
  0, 0, 0, 0,
  2.223921e-014, 3.974395e-014, 1.515518e-011, 3.254389e-011,
  0, 0, 0, 0,
  9.301416e-015, 4.14441e-014, 1.131535e-011, 2.761135e-011,
  0, 0, 0, 0,
  1.00551e-014, 4.38137e-014, 1.920455e-011, 4.099669e-011,
  0, 0, 0, 0,
  1.953908e-014, 4.993638e-014, 2.756263e-011, 5.545507e-011,
  0, 0, 0, 0,
  2.342553e-014, 7.080504e-014, 3.171327e-011, 6.462692e-011,
  0, 0, 0, 0,
  8.825192e-014, 4.507614e-014, 6.729447e-011, 1.247628e-010,
  0, 0, 0, 0,
  1.779962e-014, 5.099729e-014, 2.312783e-011, 4.264426e-011,
  0, 0, 0, 0,
  3.801007e-014, 7.792358e-014, 1.934963e-011, 4.694129e-011,
  0, 0, 0, 0,
  6.733342e-014, 1.304184e-013, 5.045298e-011, 8.488075e-011,
  0, 0, 0, 0,
  8.863635e-014, 1.242228e-013, 4.888188e-011, 8.399947e-011,
  0, 0, 0, 0,
  9.454845e-014, 1.298777e-013, 5.149978e-011, 1.060692e-010,
  0, 0, 0, 0,
  1.199243e-013, 1.412718e-013, 5.12494e-011, 1.008237e-010,
  0, 0, 0, 0,
  2.187728e-013, 1.131037e-013, 1.177371e-010, 2.093442e-010,
  0, 0, 0, 0,
  2.678623e-013, 1.524843e-013, 1.43578e-010, 2.499291e-010,
  0, 0, 0, 0,
  1.357612e-013, 8.294963e-014, 7.326899e-011, 1.25515e-010,
  0, 0, 0, 0,
  1.77574e-013, 4.984124e-014, 9.399841e-011, 1.647087e-010,
  0, 0, 0, 0,
  1.286322e-013, 6.022563e-014, 7.513862e-011, 1.403496e-010,
  0, 0, 0, 0,
  1.707957e-013, 1.023718e-013, 7.537158e-011, 1.298389e-010,
  0, 0, 0, 0,
  1.212553e-013, 5.955062e-014, 7.418362e-011, 1.309203e-010,
  0, 0, 0, 0,
  1.065059e-013, 9.421479e-014, 9.76689e-011, 1.665785e-010,
  0, 0, 0, 0,
  1.097882e-013, 1.176842e-013, 6.269999e-011, 1.155811e-010,
  0, 0, 0, 0,
  1.323992e-013, 4.135773e-014, 8.033701e-011, 1.346757e-010,
  0, 0, 0, 0,
  1.396404e-013, 4.725993e-014, 4.438558e-011, 9.261007e-011,
  0, 0, 0, 0,
  1.120939e-013, 4.687852e-014, 5.496289e-011, 1.186868e-010,
  0, 0, 0, 0,
  6.180955e-014, 4.398522e-014, 2.283523e-011, 3.675163e-011,
  0, 0, 0, 0,
  6.174236e-014, 5.496969e-014, 2.332896e-011, 4.441562e-011,
  0, 0, 0, 0,
  8.713343e-014, 4.557813e-014, 3.034589e-011, 5.00585e-011,
  0, 0, 0, 0,
  5.021734e-014, 4.241222e-014, 2.930313e-011, 4.623213e-011,
  0, 0, 0, 0,
  4.015531e-014, 1.037746e-014, 2.323519e-011, 4.160651e-011,
  0, 0, 0, 0,
  3.868536e-014, 1.389415e-014, 2.509517e-011, 4.170523e-011,
  0, 0, 0, 0,
  2.661323e-014, 1.215544e-014, 1.635883e-011, 2.811261e-011,
  0, 0, 0, 0,
  2.512915e-014, 1.830825e-014, 1.871955e-011, 3.26849e-011,
  0, 0, 0, 0,
  8.398676e-015, 1.395572e-014, 7.919924e-012, 1.471213e-011,
  0, 0, 0, 0,
  1.409558e-014, 4.053793e-014, 9.759441e-012, 2.355232e-011,
  0, 0, 0, 0,
  5.872989e-014, 2.536103e-014, 1.097698e-011, 2.505282e-011,
  0, 0, 0, 0,
  3.195224e-014, 4.780619e-014, 2.465079e-011, 5.519959e-011,
  0, 0, 0, 0,
  2.527492e-014, 5.374975e-014, 2.950523e-011, 5.819865e-011,
  0, 0, 0, 0,
  4.309769e-014, 3.394939e-014, 2.25488e-011, 4.422233e-011,
  0, 0, 0, 0,
  4.86564e-014, 3.657778e-014, 3.20059e-011, 5.707156e-011,
  0, 0, 0, 0,
  7.646376e-014, 5.165935e-014, 2.637264e-011, 5.949762e-011,
  0, 0, 0, 0,
  7.763621e-014, 3.399299e-014, 4.953723e-011, 9.714458e-011,
  0, 0, 0, 0,
  1.633705e-013, 4.579188e-014, 9.019017e-011, 1.755555e-010,
  0, 0, 0, 0,
  1.466129e-013, 4.092262e-014, 6.549412e-011, 1.193408e-010,
  0, 0, 0, 0,
  1.541867e-013, 8.57808e-014, 5.962192e-011, 1.089544e-010,
  0, 0, 0, 0,
  1.477782e-013, 3.653874e-014, 1.064955e-010, 1.860897e-010,
  0, 0, 0, 0,
  1.56098e-013, 2.676558e-014, 8.209453e-011, 1.380431e-010,
  0, 0, 0, 0,
  1.629364e-013, 4.006182e-014, 7.199031e-011, 1.223776e-010,
  0, 0, 0, 0,
  2.086666e-013, 4.420148e-014, 7.140024e-011, 1.311064e-010,
  0, 0, 0, 0,
  1.741577e-013, 4.787329e-014, 6.832737e-011, 1.341497e-010,
  0, 0, 0, 0,
  1.927033e-013, 8.038869e-014, 1.239764e-010, 2.176003e-010,
  0, 0, 0, 0,
  1.786035e-013, 6.169099e-014, 1.110316e-010, 2.031836e-010,
  0, 0, 0, 0,
  2.419244e-013, 1.070971e-013, 1.593537e-010, 2.86724e-010,
  0, 0, 0, 0,
  1.663185e-013, 1.040705e-013, 8.906615e-011, 1.83589e-010,
  0, 0, 0, 0,
  2.253494e-013, 1.062739e-013, 9.528569e-011, 1.918744e-010,
  0, 0, 0, 0,
  1.709753e-013, 8.479178e-014, 7.967951e-011, 1.335577e-010,
  0, 0, 0, 0,
  2.094137e-013, 1.227696e-013, 1.582503e-010, 2.577099e-010,
  0, 0, 0, 0,
  1.44447e-013, 7.91842e-014, 7.31064e-011, 1.286072e-010,
  0, 0, 0, 0,
  1.198197e-013, 3.695741e-014, 7.371471e-011, 1.212341e-010,
  0, 0, 0, 0,
  8.591622e-014, 3.20564e-014, 4.210406e-011, 7.415681e-011,
  0, 0, 0, 0,
  1.098951e-013, 3.721621e-014, 3.799674e-011, 7.743618e-011,
  0, 0, 0, 0,
  1.080061e-013, 3.345285e-014, 4.160365e-011, 6.88173e-011,
  0, 0, 0, 0,
  9.474945e-014, 3.537506e-014, 4.678877e-011, 8.07534e-011,
  0, 0, 0, 0,
  5.146638e-014, 2.43862e-014, 3.826996e-011, 6.929532e-011,
  0, 0, 0, 0,
  8.234574e-014, 4.730987e-014, 4.188566e-011, 8.109189e-011,
  0, 0, 0, 0,
  9.438477e-014, 2.651193e-014, 2.981411e-011, 4.864567e-011,
  0, 0, 0, 0,
  4.464607e-014, 2.575007e-014, 3.159468e-011, 5.473388e-011,
  0, 0, 0, 0,
  7.977179e-014, 4.311842e-014, 4.84454e-011, 1.02196e-010,
  0, 0, 0, 0,
  1.073313e-013, 9.879204e-014, 5.373877e-011, 1.125796e-010,
  0, 0, 0, 0,
  1.12982e-013, 7.307077e-014, 6.668151e-011, 1.106228e-010,
  0, 0, 0, 0,
  1.577534e-013, 6.487171e-014, 4.627492e-011, 8.873484e-011,
  0, 0, 0, 0,
  1.535603e-013, 8.513536e-014, 6.617918e-011, 1.17313e-010,
  0, 0, 0, 0,
  9.2545e-014, 6.382895e-014, 8.602207e-011, 1.569743e-010,
  0, 0, 0, 0,
  1.202696e-013, 6.728458e-014, 9.315946e-011, 1.59463e-010,
  0, 0, 0, 0,
  1.689864e-013, 6.991366e-014, 6.278466e-011, 1.316652e-010,
  0, 0, 0, 0,
  1.938404e-013, 6.471887e-014, 9.016056e-011, 1.637966e-010,
  0, 0, 0, 0,
  1.956319e-013, 6.488655e-014, 8.849085e-011, 1.385761e-010,
  0, 0, 0, 0,
  1.878735e-013, 6.896487e-014, 4.994753e-011, 8.289727e-011,
  0, 0, 0, 0,
  1.154254e-013, 6.565352e-014, 5.818248e-011, 1.241742e-010,
  0, 0, 0, 0,
  1.798478e-013, 5.340177e-014, 9.406273e-011, 1.71006e-010,
  0, 0, 0, 0,
  1.111811e-013, 5.885795e-014, 5.074589e-011, 9.195686e-011,
  0, 0, 0, 0,
  1.149716e-013, 5.866036e-014, 8.875272e-011, 1.752556e-010,
  0, 0, 0, 0,
  8.481977e-014, 7.247649e-014, 3.351916e-011, 6.047796e-011,
  0, 0, 0, 0,
  4.620345e-014, 6.30755e-014, 3.592278e-011, 6.084028e-011,
  0, 0, 0, 0,
  4.03432e-014, 4.992946e-014, 2.909977e-011, 6.044332e-011,
  0, 0, 0, 0,
  1.127554e-013, 8.268316e-014, 6.393708e-011, 1.157582e-010,
  0, 0, 0, 0,
  8.491912e-014, 6.308026e-014, 3.25062e-011, 5.643024e-011,
  0, 0, 0, 0,
  8.874473e-014, 6.594037e-014, 5.212466e-011, 8.633189e-011,
  0, 0, 0, 0,
  2.195838e-013, 5.554612e-014, 1.112843e-010, 1.978736e-010,
  0, 0, 0, 0,
  1.399215e-013, 6.34964e-014, 4.820966e-011, 8.529989e-011,
  0, 0, 0, 0,
  1.873267e-013, 4.936871e-014, 9.054481e-011, 1.592988e-010,
  0, 0, 0, 0,
  1.86549e-013, 7.091546e-014, 9.243958e-011, 1.576652e-010,
  0, 0, 0, 0,
  1.627911e-013, 1.112453e-013, 1.131933e-010, 2.012893e-010,
  0, 0, 0, 0,
  2.676761e-013, 7.805974e-014, 1.145421e-010, 2.233239e-010,
  0, 0, 0, 0,
  2.077441e-013, 8.672918e-014, 9.662943e-011, 1.75796e-010,
  0, 0, 0, 0,
  2.050307e-013, 1.023845e-013, 1.314537e-010, 2.212227e-010,
  0, 0, 0, 0,
  1.905602e-013, 7.71628e-014, 1.121969e-010, 1.947952e-010,
  0, 0, 0, 0,
  2.279364e-013, 1.019524e-013, 1.255321e-010, 2.096798e-010,
  0, 0, 0, 0,
  1.592806e-013, 9.639526e-014, 7.719238e-011, 1.350338e-010,
  0, 0, 0, 0,
  1.865122e-013, 5.846259e-014, 7.952285e-011, 1.515984e-010,
  0, 0, 0, 0,
  1.574207e-013, 6.165666e-014, 7.249199e-011, 1.372154e-010,
  0, 0, 0, 0,
  1.332662e-013, 4.528443e-014, 5.106742e-011, 1.081022e-010,
  0, 0, 0, 0,
  1.613148e-013, 6.087717e-014, 4.149878e-011, 5.800142e-011,
  0, 0, 0, 0,
  8.35666e-014, 9.478261e-014, 5.681178e-011, 1.045332e-010,
  0, 0, 0, 0,
  1.560558e-013, 5.587175e-014, 8.967939e-011, 1.632946e-010,
  0, 0, 0, 0,
  1.028884e-013, 7.017402e-014, 5.033851e-011, 9.735228e-011,
  0, 0, 0, 0,
  1.292633e-013, 7.998695e-014, 5.092635e-011, 7.957107e-011,
  0, 0, 0, 0,
  1.838518e-013, 8.425878e-014, 7.602707e-011, 1.309168e-010,
  0, 0, 0, 0,
  1.60604e-013, 6.809318e-014, 9.220167e-011, 1.417118e-010,
  0, 0, 0, 0,
  1.022825e-013, 5.649902e-014, 6.129926e-011, 1.119598e-010,
  0, 0, 0, 0,
  1.390292e-013, 4.723888e-014, 6.666395e-011, 1.117008e-010,
  0, 0, 0, 0,
  1.393796e-013, 6.689953e-014, 7.88736e-011, 1.518891e-010,
  0, 0, 0, 0,
  2.115105e-013, 9.090219e-014, 7.916579e-011, 1.289742e-010,
  0, 0, 0, 0,
  1.548877e-013, 8.27085e-014, 7.302323e-011, 1.290894e-010,
  0, 0, 0, 0,
  2.145585e-013, 8.541118e-014, 7.281686e-011, 1.20892e-010,
  0, 0, 0, 0,
  2.387194e-013, 1.234511e-013, 1.206106e-010, 2.362039e-010,
  0, 0, 0, 0,
  2.30924e-013, 9.026924e-014, 1.31117e-010, 2.296299e-010,
  0, 0, 0, 0,
  1.387223e-013, 1.441122e-013, 7.864052e-011, 1.30972e-010,
  0, 0, 0, 0,
  2.204804e-013, 1.391864e-013, 1.701096e-010, 3.115944e-010,
  0, 0, 0, 0,
  1.64825e-013, 9.750219e-014, 1.08695e-010, 2.069813e-010,
  0, 0, 0, 0,
  5.515654e-015, 3.592953e-015, 2.8598e-012, 4.403021e-012,
  0, 0, 0, 0,
  3.135077e-014, 5.642602e-015, 3.177905e-011, 2.660486e-011,
  0, 0, 0, 0,
  1.063629e-013, 1.684421e-014, 5.253637e-012, 4.279432e-012,
  0, 0, 0, 0,
  1.213437e-014, 1.697871e-014, 9.905288e-012, 1.472136e-011,
  0, 0, 0, 0,
  7.474464e-015, 5.273974e-015, 3.590521e-012, 4.628406e-012,
  0, 0, 0, 0,
  5.783799e-015, 2.556109e-015, 1.313439e-011, 1.343565e-011,
  0, 0, 0, 0,
  8.706145e-014, 1.663938e-014, 1.048865e-011, 9.748722e-012,
  0, 0, 0, 0,
  3.426983e-015, 1.515395e-014, 8.939348e-012, 1.890922e-011,
  0, 0, 0, 0,
  4.57351e-015, 3.587648e-015, 1.859393e-011, 9.415954e-012,
  0, 0, 0, 0,
  3.117866e-014, 2.016009e-013, 1.644429e-011, 1.082141e-011,
  0, 0, 0, 0,
  8.506805e-014, 1.574771e-014, 2.850316e-012, 2.987845e-012,
  0, 0, 0, 0,
  1.029156e-014, 2.887489e-015, 2.853783e-012, 3.085533e-012,
  0, 0, 0, 0,
  2.312475e-015, 3.780243e-015, 7.090996e-012, 8.524361e-012,
  0, 0, 0, 0,
  4.505029e-015, 2.709038e-015, 4.066261e-012, 4.394381e-012,
  0, 0, 0, 0,
  2.997411e-015, 1.922892e-015, 2.704505e-012, 2.721859e-012,
  0, 0, 0, 0,
  3.884921e-015, 2.857802e-015, 4.329349e-012, 6.006906e-012,
  0, 0, 0, 0,
  8.170529e-015, 2.365194e-015, 7.331742e-012, 1.234399e-011,
  0, 0, 0, 0,
  2.274914e-015, 3.374481e-015, 2.802279e-012, 4.2164e-012,
  0, 0, 0, 0,
  3.266185e-015, 1.404299e-014, 2.787437e-012, 3.888156e-012,
  0, 0, 0, 0,
  3.644583e-015, 6.329542e-015, 5.71528e-012, 1.174206e-011,
  0, 0, 0, 0,
  2.567177e-015, 2.534422e-015, 5.040586e-012, 9.638674e-012,
  0, 0, 0, 0,
  3.020717e-015, 3.21763e-015, 3.200669e-012, 4.16478e-012,
  0, 0, 0, 0,
  1.130998e-014, 3.717882e-015, 5.345218e-012, 8.647945e-012,
  0, 0, 0, 0,
  8.622103e-014, 1.372731e-014, 8.486926e-012, 1.172655e-011,
  0, 0, 0, 0,
  2.470357e-015, 1.091509e-014, 7.23741e-012, 1.029633e-011,
  0, 0, 0, 0,
  2.660227e-015, 6.646409e-015, 8.179148e-012, 8.672773e-012,
  0, 0, 0, 0,
  5.227925e-015, 8.432674e-015, 4.454238e-012, 7.911816e-012,
  0, 0, 0, 0,
  9.382834e-014, 1.530867e-014, 1.252481e-011, 1.509205e-011,
  0, 0, 0, 0,
  5.154983e-015, 7.183974e-015, 3.637937e-012, 6.585656e-012,
  0, 0, 0, 0,
  4.019997e-015, 2.412945e-015, 6.124531e-012, 7.229317e-012,
  0, 0, 0, 0,
  3.005524e-015, 3.374573e-015, 3.587844e-012, 1.803573e-012,
  0, 0, 0, 0,
  3.399553e-015, 3.964253e-015, 5.741279e-012, 8.86603e-012,
  0, 0, 0, 0,
  3.109508e-015, 2.859076e-015, 3.005131e-012, 4.426971e-012,
  0, 0, 0, 0,
  1.128388e-014, 3.004297e-015, 4.352751e-012, 1.570117e-011,
  0, 0, 0, 0,
  5.573246e-015, 3.006603e-015, 6.223163e-012, 9.849546e-012,
  0, 0, 0, 0,
  7.199207e-014, 1.162831e-014, 4.828566e-012, 6.501555e-012,
  0, 0, 0, 0,
  8.570705e-014, 1.34303e-014, 1.166732e-011, 2.207039e-011,
  0, 0, 0, 0,
  3.117586e-015, 3.601329e-015, 3.510643e-012, 5.150168e-012,
  0, 0, 0, 0,
  6.678078e-015, 2.901463e-015, 2.010043e-012, 1.651926e-012,
  0, 0, 0, 0,
  1.499963e-014, 3.567314e-015, 2.276193e-012, 3.110054e-012,
  0, 0, 0, 0,
  7.596734e-014, 1.203306e-014, 3.498653e-012, 3.50681e-012,
  0, 0, 0, 0,
  5.347533e-015, 3.459049e-015, 5.60039e-012, 8.426817e-012,
  0, 0, 0, 0,
  3.134097e-015, 3.146343e-015, 3.58079e-012, 5.539821e-012,
  0, 0, 0, 0,
  3.540537e-015, 1.927372e-015, 3.311687e-012, 4.042816e-012,
  0, 0, 0, 0,
  9.19902e-014, 1.434918e-014, 2.65749e-012, 2.420461e-012,
  0, 0, 0, 0,
  9.037892e-015, 5.24283e-015, 3.453028e-012, 5.185845e-012,
  0, 0, 0, 0,
  4.490575e-015, 2.113497e-014, 5.154493e-012, 1.223758e-011,
  0, 0, 0, 0,
  4.342363e-015, 1.001523e-014, 3.134059e-012, 3.104224e-012,
  0, 0, 0, 0,
  1.285033e-013, 5.487652e-014, 7.38131e-012, 1.705171e-011,
  0, 0, 0, 0,
  1.81868e-014, 4.855956e-015, 1.61478e-011, 2.113551e-011,
  0, 0, 0, 0,
  2.698958e-015, 3.580984e-015, 2.928759e-012, 2.727108e-012,
  0, 0, 0, 0,
  2.147343e-015, 2.271856e-015, 2.051061e-012, 1.650367e-012,
  0, 0, 0, 0,
  4.670792e-014, 8.557807e-015, 2.90252e-012, 3.663896e-012,
  0, 0, 0, 0,
  3.657848e-014, 6.541995e-015, 3.814836e-012, 6.770717e-012,
  0, 0, 0, 0,
  2.292725e-015, 2.29745e-015, 2.826823e-012, 2.560904e-012,
  0, 0, 0, 0,
  3.228907e-015, 3.112696e-015, 2.51065e-012, 2.064431e-012,
  0, 0, 0, 0,
  2.567494e-014, 5.609828e-015, 1.796171e-012, 2.112094e-012,
  0, 0, 0, 0,
  6.490143e-014, 1.079736e-014, 3.521714e-012, 3.406107e-012,
  0, 0, 0, 0,
  3.714051e-015, 4.454221e-015, 2.141554e-012, 3.180296e-012,
  0, 0, 0, 0,
  2.042274e-015, 2.89254e-015, 1.005027e-012, 1.960574e-012,
  0, 0, 0, 0,
  3.616576e-015, 2.364425e-015, 2.337638e-012, 2.51174e-012,
  0, 0, 0, 0,
  1.774858e-015, 2.35431e-015, 1.899469e-012, 2.097493e-012,
  0, 0, 0, 0,
  3.209478e-015, 2.70567e-015, 2.786889e-012, 2.621247e-012,
  0, 0, 0, 0,
  2.23519e-015, 2.624824e-015, 1.452104e-012, 1.568284e-012,
  0, 0, 0, 0,
  3.796239e-015, 3.281407e-015, 2.452827e-012, 2.080343e-012,
  0, 0, 0, 0,
  1.317498e-013, 2.312249e-014, 3.751438e-012, 6.414667e-012,
  0, 0, 0, 0,
  4.971295e-015, 5.603871e-015, 3.092899e-012, 4.306609e-012,
  0, 0, 0, 0,
  5.603527e-015, 2.405912e-014, 1.443233e-011, 2.64208e-011,
  0, 0, 0, 0,
  5.213611e-015, 2.190532e-014, 1.512917e-011, 2.619814e-011,
  0, 0, 0, 0,
  6.758948e-014, 1.154927e-014, 3.468219e-012, 7.040177e-012,
  0, 0, 0, 0,
  1.967296e-014, 4.081532e-015, 2.476785e-012, 2.78484e-012,
  0, 0, 0, 0,
  7.520939e-015, 4.736126e-015, 1.312118e-011, 1.357028e-011,
  0, 0, 0, 0,
  5.075633e-015, 3.132247e-015, 2.518746e-012, 3.476838e-012,
  0, 0, 0, 0,
  3.765619e-014, 6.70758e-015, 2.047118e-012, 2.409311e-012,
  0, 0, 0, 0,
  5.280418e-014, 8.605247e-015, 2.300944e-012, 2.288001e-012,
  0, 0, 0, 0,
  4.056312e-015, 2.334647e-015, 2.675645e-012, 2.4023e-012,
  0, 0, 0, 0,
  6.259946e-015, 2.966516e-015, 1.877946e-012, 2.070817e-012,
  0, 0, 0, 0,
  8.830534e-015, 3.358418e-015, 6.682193e-012, 9.025461e-012,
  0, 0, 0, 0,
  9.021468e-015, 4.565818e-015, 9.835322e-012, 1.390456e-011,
  0, 0, 0, 0,
  7.293414e-015, 7.247828e-015, 4.954758e-012, 9.465886e-012,
  0, 0, 0, 0,
  5.759351e-015, 5.292277e-015, 7.399052e-012, 8.043131e-012,
  0, 0, 0, 0,
  6.466452e-015, 9.586207e-015, 8.681395e-012, 1.487487e-011,
  0, 0, 0, 0,
  1.39388e-013, 2.224751e-014, 6.200661e-012, 9.522955e-012,
  0, 0, 0, 0,
  7.445025e-015, 1.281736e-014, 8.030379e-012, 1.509475e-011,
  0, 0, 0, 0,
  5.665572e-015, 7.907752e-015, 6.989156e-012, 1.224051e-011,
  0, 0, 0, 0,
  3.910986e-015, 5.641056e-015, 6.351818e-012, 8.61884e-012,
  0, 0, 0, 0,
  7.610561e-014, 1.274844e-014, 5.186936e-012, 6.969697e-012,
  0, 0, 0, 0,
  1.1814e-014, 1.072012e-014, 6.001407e-012, 1.106861e-011,
  0, 0, 0, 0,
  5.778743e-015, 5.91348e-015, 4.488845e-012, 7.308779e-012,
  0, 0, 0, 0,
  5.815249e-015, 3.11975e-014, 1.583078e-011, 2.762631e-011,
  0, 0, 0, 0,
  5.770577e-014, 2.102443e-014, 1.386889e-011, 2.250035e-011,
  0, 0, 0, 0,
  3.439056e-014, 1.084296e-014, 8.344361e-012, 1.461035e-011,
  0, 0, 0, 0,
  7.375094e-015, 1.766425e-014, 1.231553e-011, 2.494825e-011,
  0, 0, 0, 0,
  1.309975e-014, 5.40622e-015, 1.504445e-011, 1.678487e-011,
  0, 0, 0, 0,
  1.6978e-014, 1.335854e-014, 1.169331e-011, 2.582981e-011,
  0, 0, 0, 0,
  3.376234e-015, 4.568567e-015, 5.485017e-012, 6.582252e-012,
  0, 0, 0, 0,
  4.064147e-015, 3.558005e-015, 2.627427e-012, 5.123948e-012,
  0, 0, 0, 0,
  3.64619e-015, 4.452091e-015, 4.127126e-012, 4.473302e-012,
  0, 0, 0, 0,
  5.651686e-015, 4.059077e-015, 3.492242e-012, 3.956699e-012,
  0, 0, 0, 0,
  5.891139e-015, 2.841249e-015, 3.017936e-012, 2.703833e-012,
  0, 0, 0, 0,
  3.233431e-015, 5.196139e-015, 2.015673e-012, 1.858436e-012,
  0, 0, 0, 0,
  7.383059e-015, 3.862348e-014, 2.035718e-012, 1.97751e-012,
  0, 0, 0, 0,
  9.187142e-014, 1.573971e-014, 1.348957e-011, 2.81138e-011,
  0, 0, 0, 0,
  3.265522e-014, 6.993165e-015, 5.242329e-011, 6.295167e-011,
  0, 0, 0, 0,
  1.209842e-014, 1.066931e-014, 5.482705e-011, 5.561637e-011,
  0, 0, 0, 0,
  7.024152e-014, 2.711328e-014, 2.334766e-011, 6.113415e-011,
  0, 0, 0, 0,
  5.729629e-015, 5.898385e-015, 4.817139e-012, 8.163348e-012,
  0, 0, 0, 0,
  8.529408e-015, 9.686451e-015, 6.22156e-012, 1.218883e-011,
  0, 0, 0, 0,
  2.419905e-014, 1.334203e-014, 3.136367e-011, 6.372021e-011,
  0, 0, 0, 0,
  1.492896e-014, 5.126055e-015, 3.728849e-012, 7.940785e-012,
  0, 0, 0, 0,
  1.052894e-014, 4.931647e-015, 5.341538e-012, 7.45639e-012,
  0, 0, 0, 0,
  1.711364e-014, 4.255395e-015, 2.230803e-012, 7.183662e-012,
  0, 0, 0, 0,
  1.368361e-014, 6.800944e-015, 2.827912e-012, 7.88973e-012,
  0, 0, 0, 0,
  3.134021e-014, 7.196846e-015, 4.245844e-012, 1.258658e-011,
  0, 0, 0, 0,
  5.539834e-014, 1.041951e-014, 7.608632e-012, 2.234564e-011,
  0, 0, 0, 0,
  4.694209e-014, 9.967428e-015, 1.872218e-011, 3.585736e-011,
  0, 0, 0, 0,
  5.1889e-014, 1.135223e-014, 4.47223e-012, 1.259959e-011,
  0, 0, 0, 0,
  5.488958e-014, 1.89367e-014, 4.256926e-012, 8.935968e-012,
  0, 0, 0, 0,
  1.676843e-013, 3.484568e-014, 6.280693e-012, 2.984671e-011,
  0, 0, 0, 0,
  4.581993e-013, 7.552326e-014, 9.929274e-012, 5.032648e-011,
  0, 0, 0, 0,
  3.399251e-013, 6.685592e-014, 7.030674e-012, 3.592591e-011,
  0, 0, 0, 0,
  6.93033e-013, 1.287553e-013, 2.24226e-011, 9.075114e-011,
  0, 0, 0, 0,
  5.768942e-013, 1.283378e-013, 1.517396e-011, 5.82682e-011,
  0, 0, 0, 0,
  1.432512e-012, 2.991457e-013, 4.922088e-011, 2.109205e-010,
  0, 0, 0, 0,
  2.461783e-012, 4.888683e-013, 1.383483e-010, 4.633711e-010,
  0, 0, 0, 0,
  2.047318e-012, 6.298118e-013, 9.609138e-011, 3.465039e-010,
  0, 0, 0, 0,
  3.555091e-012, 1.133918e-012, 1.748902e-010, 6.732134e-010,
  0, 0, 0, 0,
  9.052324e-012, 2.492426e-012, 7.168341e-010, 2.075758e-009,
  0, 0, 0, 0,
  1.576668e-011, 4.597327e-012, 1.452827e-009, 7.355372e-009,
  0, 0, 0, 0,
  2.312177e-011, 5.907883e-012, 1.367543e-009, 5.269294e-009,
  0, 0, 0, 0,
  1.210831e-011, 4.066984e-012, 9.899134e-010, 3.386681e-009,
  0, 0, 0, 0,
  1.854973e-011, 5.696314e-012, 1.303788e-009, 4.501334e-009,
  0, 0, 0, 0,
  1.587141e-011, 6.40848e-012, 1.354473e-009, 5.44145e-009,
  0, 0, 0, 0,
  5.473583e-012, 2.251197e-012, 4.04225e-010, 1.702232e-009,
  0, 0, 0, 0,
  3.798028e-012, 8.688161e-013, 1.485468e-010, 6.526484e-010,
  0, 0, 0, 0,
  2.429548e-012, 5.034493e-013, 8.122103e-011, 3.564427e-010,
  0, 0, 0, 0,
  1.977008e-012, 5.033163e-013, 6.99435e-011, 3.071345e-010,
  0, 0, 0, 0,
  8.831093e-013, 3.48226e-013, 5.920268e-011, 1.766047e-010,
  0, 0, 0, 0,
  5.575158e-013, 2.81877e-013, 5.006727e-011, 1.521321e-010,
  0, 0, 0, 0,
  3.177486e-013, 2.599423e-013, 2.488272e-011, 7.797949e-011,
  0, 0, 0, 0,
  4.928655e-013, 2.259247e-013, 2.329966e-011, 6.144919e-011,
  0, 0, 0, 0,
  3.259296e-013, 9.150593e-014, 1.694059e-011, 5.34545e-011,
  0, 0, 0, 0,
  3.021177e-013, 6.00953e-014, 1.544644e-011, 4.120956e-011,
  0, 0, 0, 0,
  8.415713e-014, 2.819586e-014, 8.644361e-012, 2.022831e-011,
  0, 0, 0, 0,
  1.256387e-013, 2.900514e-014, 9.824372e-012, 3.120537e-011,
  0, 0, 0, 0,
  5.23532e-014, 1.220057e-013, 6.101802e-011, 1.450683e-010,
  0, 0, 0, 0,
  3.143081e-014, 2.0496e-014, 9.892397e-012, 1.926832e-011,
  0, 0, 0, 0,
  2.201717e-014, 2.451992e-014, 9.847022e-012, 2.228489e-011,
  0, 0, 0, 0,
  1.486505e-014, 1.70148e-014, 1.367693e-011, 2.937734e-011,
  0, 0, 0, 0,
  2.34352e-014, 2.458283e-014, 1.365358e-011, 2.508365e-011,
  0, 0, 0, 0,
  2.185204e-014, 1.010722e-013, 5.057255e-011, 1.194404e-010,
  0, 0, 0, 0,
  3.333672e-014, 7.975734e-014, 4.723734e-011, 1.025383e-010,
  0, 0, 0, 0,
  2.351056e-014, 7.924941e-014, 4.983764e-011, 1.217851e-010,
  0, 0, 0, 0,
  7.81714e-014, 9.142011e-014, 3.473752e-011, 7.047441e-011,
  0, 0, 0, 0,
  1.513718e-014, 7.398862e-014, 2.941106e-011, 6.544374e-011,
  0, 0, 0, 0,
  1.686504e-014, 9.836054e-014, 4.612007e-011, 1.060056e-010,
  0, 0, 0, 0,
  8.665918e-015, 3.103273e-014, 1.620968e-011, 3.286379e-011,
  0, 0, 0, 0,
  6.527328e-015, 3.641512e-014, 1.705473e-011, 4.078534e-011,
  0, 0, 0, 0,
  7.586911e-015, 3.540422e-014, 2.11522e-011, 5.068044e-011,
  0, 0, 0, 0,
  6.646351e-015, 1.352548e-014, 1.201397e-011, 1.413372e-011,
  0, 0, 0, 0,
  4.002493e-015, 9.648186e-015, 7.72327e-012, 1.528986e-011,
  0, 0, 0, 0,
  5.127713e-015, 2.744882e-014, 1.607946e-011, 3.715086e-011,
  0, 0, 0, 0,
  4.586098e-015, 1.338668e-014, 7.530711e-012, 1.480617e-011,
  0, 0, 0, 0,
  6.024676e-015, 1.038776e-014, 6.938447e-012, 1.205057e-011,
  0, 0, 0, 0,
  3.700634e-015, 1.462195e-014, 6.455648e-012, 1.599645e-011,
  0, 0, 0, 0,
  1.950137e-014, 3.264782e-014, 1.657273e-011, 4.040209e-011,
  0, 0, 0, 0,
  4.973882e-015, 2.161083e-014, 1.088946e-011, 2.309425e-011,
  0, 0, 0, 0,
  8.81249e-015, 4.865195e-014, 2.932379e-011, 6.607751e-011,
  0, 0, 0, 0,
  1.26917e-014, 7.086916e-014, 3.421088e-011, 9.237296e-011,
  0, 0, 0, 0,
  3.450267e-014, 1.998027e-013, 5.703614e-011, 1.527425e-010,
  0, 0, 0, 0,
  1.314437e-013, 6.739357e-014, 2.542613e-011, 6.008267e-011,
  0, 0, 0, 0,
  2.421454e-014, 1.499363e-013, 4.415314e-011, 1.00713e-010,
  0, 0, 0, 0,
  2.167917e-014, 9.638917e-014, 3.211336e-011, 8.700771e-011,
  0, 0, 0, 0,
  1.060273e-014, 4.399491e-014, 2.267316e-011, 5.381098e-011,
  0, 0, 0, 0,
  7.369627e-014, 5.221546e-014, 1.579632e-011, 3.959264e-011,
  0, 0, 0, 0,
  1.405002e-014, 4.373379e-014, 2.177748e-011, 5.27208e-011,
  0, 0, 0, 0,
  5.80993e-015, 2.988415e-014, 1.532539e-011, 3.580162e-011,
  0, 0, 0, 0,
  7.995966e-015, 4.22677e-014, 1.432116e-011, 3.500687e-011,
  0, 0, 0, 0,
  5.452046e-014, 6.018502e-014, 3.776109e-011, 8.99003e-011,
  0, 0, 0, 0,
  3.460877e-014, 3.820903e-014, 2.536253e-011, 5.545581e-011,
  0, 0, 0, 0,
  1.631065e-014, 7.112368e-014, 4.547351e-011, 9.599912e-011,
  0, 0, 0, 0,
  1.288045e-014, 5.009363e-014, 2.63227e-011, 6.233495e-011,
  0, 0, 0, 0,
  1.241632e-014, 4.060064e-014, 3.025614e-011, 7.04774e-011,
  0, 0, 0, 0,
  1.638138e-014, 3.559043e-014, 2.581501e-011, 5.208509e-011,
  0, 0, 0, 0,
  1.241566e-014, 6.453549e-014, 5.091648e-011, 1.183531e-010,
  0, 0, 0, 0,
  1.061188e-014, 5.648017e-014, 2.963751e-011, 6.81721e-011,
  0, 0, 0, 0,
  1.902039e-014, 1.172668e-013, 3.938302e-011, 7.811214e-011,
  0, 0, 0, 0,
  1.287397e-013, 5.562834e-014, 2.895113e-011, 6.762663e-011,
  0, 0, 0, 0,
  2.054362e-014, 1.121353e-013, 5.917201e-011, 1.387041e-010,
  0, 0, 0, 0,
  1.332293e-014, 7.073624e-014, 3.952154e-011, 9.356745e-011,
  0, 0, 0, 0,
  1.301282e-014, 8.093493e-014, 3.604719e-011, 8.861306e-011,
  0, 0, 0, 0,
  7.90197e-014, 2.11705e-014, 1.072897e-011, 2.142408e-011,
  0, 0, 0, 0,
  7.159682e-015, 2.022056e-014, 1.794761e-011, 3.372721e-011,
  0, 0, 0, 0,
  1.125707e-014, 6.888557e-014, 3.251723e-011, 7.688431e-011,
  0, 0, 0, 0,
  8.654812e-015, 4.228675e-014, 1.80911e-011, 4.706882e-011,
  0, 0, 0, 0,
  6.392434e-014, 1.758306e-014, 1.119037e-011, 1.909465e-011,
  0, 0, 0, 0,
  2.264865e-014, 1.094123e-014, 7.735592e-012, 1.333575e-011,
  0, 0, 0, 0,
  3.211111e-015, 1.24099e-014, 5.667794e-012, 1.502579e-011,
  0, 0, 0, 0,
  4.529109e-015, 1.140369e-014, 8.794771e-012, 1.901035e-011,
  0, 0, 0, 0,
  6.535492e-015, 3.010054e-014, 1.837368e-011, 3.957294e-011,
  0, 0, 0, 0,
  6.912887e-015, 4.064834e-014, 2.331914e-011, 5.525775e-011,
  0, 0, 0, 0,
  5.758733e-015, 3.040723e-014, 1.982724e-011, 3.993683e-011,
  0, 0, 0, 0,
  8.434747e-015, 4.549171e-014, 2.671349e-011, 6.001121e-011,
  0, 0, 0, 0,
  2.212964e-014, 3.805294e-014, 1.937485e-011, 5.204506e-011,
  0, 0, 0, 0,
  1.161059e-013, 4.628049e-014, 3.896867e-011, 9.930837e-011,
  0, 0, 0, 0,
  7.538037e-015, 3.321544e-014, 1.525664e-011, 2.67292e-011,
  0, 0, 0, 0,
  2.426342e-014, 1.080761e-013, 5.515339e-011, 1.186888e-010,
  0, 0, 0, 0,
  7.162724e-014, 1.627206e-013, 8.287555e-011, 1.797221e-010,
  0, 0, 0, 0,
  7.894096e-014, 1.380334e-013, 6.160276e-011, 1.177505e-010,
  0, 0, 0, 0,
  3.822053e-014, 1.439289e-013, 5.39364e-011, 1.272429e-010,
  0, 0, 0, 0,
  7.782238e-014, 1.949978e-013, 6.113963e-011, 1.343975e-010,
  0, 0, 0, 0,
  4.533293e-014, 5.497998e-014, 6.214351e-011, 1.186467e-010,
  0, 0, 0, 0,
  7.630983e-014, 8.757924e-014, 6.189792e-011, 1.216026e-010,
  0, 0, 0, 0,
  4.303203e-014, 5.843933e-014, 4.945334e-011, 1.032063e-010,
  0, 0, 0, 0,
  9.825615e-014, 3.732016e-014, 6.999194e-011, 1.457974e-010,
  0, 0, 0, 0,
  7.9799e-014, 5.70109e-014, 4.57646e-011, 9.595353e-011,
  0, 0, 0, 0,
  1.23806e-013, 1.311757e-013, 9.333607e-011, 2.265631e-010,
  0, 0, 0, 0,
  9.077092e-014, 8.31348e-014, 4.782914e-011, 8.967566e-011,
  0, 0, 0, 0,
  1.428929e-013, 1.075902e-013, 6.894371e-011, 1.90682e-010,
  0, 0, 0, 0,
  8.809109e-014, 8.019085e-014, 5.68639e-011, 1.510107e-010,
  0, 0, 0, 0,
  4.186909e-014, 4.72645e-014, 3.668845e-011, 9.189597e-011,
  0, 0, 0, 0,
  6.701373e-014, 4.885708e-014, 2.89446e-011, 7.457001e-011,
  0, 0, 0, 0,
  1.360855e-013, 7.149435e-014, 5.332317e-011, 1.449029e-010,
  0, 0, 0, 0,
  1.755113e-014, 2.31859e-014, 2.170025e-011, 3.759861e-011,
  0, 0, 0, 0,
  1.543802e-014, 1.589394e-014, 1.655614e-011, 2.823099e-011,
  0, 0, 0, 0,
  9.435702e-014, 2.365098e-014, 1.705236e-011, 3.750414e-011,
  0, 0, 0, 0,
  1.54729e-014, 2.805506e-014, 1.805766e-011, 3.759786e-011,
  0, 0, 0, 0,
  1.159679e-014, 4.178795e-015, 7.95628e-012, 1.564408e-011,
  0, 0, 0, 0,
  1.906941e-014, 6.57841e-015, 7.608329e-012, 1.52047e-011,
  0, 0, 0, 0,
  7.213593e-015, 9.096804e-015, 7.784317e-012, 1.857571e-011,
  0, 0, 0, 0,
  8.190133e-015, 6.77905e-015, 5.284939e-012, 8.520017e-012,
  0, 0, 0, 0,
  4.004816e-015, 7.453193e-015, 6.869097e-012, 9.704446e-012,
  0, 0, 0, 0,
  1.264268e-014, 1.411173e-014, 7.625751e-012, 1.493186e-011,
  0, 0, 0, 0,
  5.741298e-014, 1.983892e-014, 1.137629e-011, 2.569057e-011,
  0, 0, 0, 0,
  2.81437e-014, 3.24292e-014, 1.989848e-011, 4.720769e-011,
  0, 0, 0, 0,
  1.239254e-014, 4.483988e-014, 1.503059e-011, 3.176905e-011,
  0, 0, 0, 0,
  7.138206e-015, 2.643997e-014, 1.996414e-011, 4.344305e-011,
  0, 0, 0, 0,
  3.128171e-014, 1.416038e-014, 1.35124e-011, 2.454226e-011,
  0, 0, 0, 0,
  6.164756e-014, 2.9702e-014, 2.398546e-011, 5.024823e-011,
  0, 0, 0, 0,
  9.032949e-014, 3.114691e-014, 1.946747e-011, 7.324883e-011,
  0, 0, 0, 0,
  7.822473e-014, 2.190354e-014, 2.54662e-011, 6.946024e-011,
  0, 0, 0, 0,
  9.258096e-014, 2.785343e-014, 4.403419e-011, 1.164661e-010,
  0, 0, 0, 0,
  2.134145e-013, 4.995027e-014, 6.583005e-011, 1.441086e-010,
  0, 0, 0, 0,
  7.019438e-014, 1.546481e-014, 3.456547e-011, 6.990606e-011,
  0, 0, 0, 0,
  5.632157e-014, 1.039942e-014, 2.442833e-011, 5.18019e-011,
  0, 0, 0, 0,
  1.579067e-013, 3.267451e-014, 5.279182e-011, 1.264405e-010,
  0, 0, 0, 0,
  3.02321e-013, 4.975329e-014, 7.70938e-011, 2.481583e-010,
  0, 0, 0, 0,
  8.101039e-014, 3.879393e-014, 7.401273e-011, 1.446717e-010,
  0, 0, 0, 0,
  1.09937e-013, 4.480243e-014, 6.706302e-011, 1.364099e-010,
  0, 0, 0, 0,
  1.424138e-013, 4.283993e-014, 6.594825e-011, 1.587512e-010,
  0, 0, 0, 0,
  2.347428e-013, 1.067449e-013, 5.898514e-011, 1.481763e-010,
  0, 0, 0, 0,
  2.324747e-013, 1.000188e-013, 6.37004e-011, 1.960331e-010,
  0, 0, 0, 0,
  1.94927e-013, 6.837261e-014, 6.200916e-011, 1.638039e-010,
  0, 0, 0, 0,
  2.044635e-013, 7.41637e-014, 8.542654e-011, 2.396752e-010,
  0, 0, 0, 0,
  6.242589e-013, 1.495225e-013, 1.951656e-010, 5.536638e-010,
  0, 0, 0, 0,
  8.431274e-014, 5.589346e-014, 5.449523e-011, 1.313027e-010,
  0, 0, 0, 0,
  3.738855e-014, 4.044548e-014, 3.958411e-011, 7.896472e-011,
  0, 0, 0, 0,
  2.441177e-014, 2.026833e-014, 2.952169e-011, 5.571998e-011,
  0, 0, 0, 0,
  8.3437e-014, 2.828783e-014, 3.02082e-011, 8.498757e-011,
  0, 0, 0, 0,
  8.641715e-014, 1.568072e-014, 1.672473e-011, 4.090652e-011,
  0, 0, 0, 0,
  3.687546e-014, 3.149865e-014, 2.559753e-011, 5.844551e-011,
  0, 0, 0, 0,
  1.425891e-014, 1.203514e-014, 1.123953e-011, 2.985025e-011,
  0, 0, 0, 0,
  1.408618e-014, 1.202764e-014, 1.752392e-011, 3.36226e-011,
  0, 0, 0, 0,
  8.676781e-014, 1.566195e-014, 1.17831e-011, 2.690185e-011,
  0, 0, 0, 0,
  1.02246e-014, 1.713784e-014, 1.133729e-011, 2.265601e-011,
  0, 0, 0, 0,
  6.32034e-014, 6.047519e-014, 4.091897e-011, 9.701867e-011,
  0, 0, 0, 0,
  6.766379e-014, 1.618496e-013, 8.831394e-011, 2.04051e-010,
  0, 0, 0, 0,
  4.861797e-014, 4.258261e-014, 4.616159e-011, 1.100096e-010,
  0, 0, 0, 0,
  3.446683e-014, 4.183377e-014, 3.215571e-011, 8.262124e-011,
  0, 0, 0, 0,
  3.881914e-014, 6.740677e-014, 3.968433e-011, 8.317191e-011,
  0, 0, 0, 0,
  1.136895e-013, 7.276626e-014, 3.436013e-011, 9.341257e-011,
  0, 0, 0, 0,
  1.400558e-013, 8.019194e-014, 7.605387e-011, 2.016244e-010,
  0, 0, 0, 0,
  1.26138e-013, 4.618972e-014, 5.473855e-011, 1.43784e-010,
  0, 0, 0, 0,
  6.850472e-014, 4.601379e-014, 4.378293e-011, 1.050426e-010,
  0, 0, 0, 0,
  4.284307e-014, 4.601097e-014, 5.122266e-011, 1.079794e-010,
  0, 0, 0, 0,
  9.303689e-014, 3.351231e-014, 4.537528e-011, 9.588022e-011,
  0, 0, 0, 0,
  1.206962e-013, 3.046688e-014, 3.621276e-011, 8.745027e-011,
  0, 0, 0, 0,
  8.33024e-014, 4.547742e-014, 5.227347e-011, 1.352088e-010,
  0, 0, 0, 0,
  3.63863e-014, 3.446978e-014, 3.229244e-011, 6.371736e-011,
  0, 0, 0, 0,
  4.177149e-014, 3.119178e-014, 2.46302e-011, 6.584563e-011,
  0, 0, 0, 0,
  8.235198e-014, 3.346685e-014, 2.698273e-011, 5.805602e-011,
  0, 0, 0, 0,
  1.590728e-014, 2.812954e-014, 3.110615e-011, 5.581639e-011,
  0, 0, 0, 0,
  3.297034e-014, 5.970873e-014, 2.127168e-011, 5.013803e-011,
  0, 0, 0, 0,
  1.457122e-013, 4.729765e-014, 5.398348e-011, 1.60947e-010,
  0, 0, 0, 0,
  6.972543e-014, 5.119768e-014, 3.346589e-011, 9.471115e-011,
  0, 0, 0, 0,
  3.009024e-014, 3.684366e-014, 2.16412e-011, 4.577903e-011,
  0, 0, 0, 0,
  4.554055e-014, 3.1018e-014, 2.826383e-011, 6.230604e-011,
  0, 0, 0, 0,
  4.668213e-014, 3.100691e-014, 2.564488e-011, 5.833754e-011,
  0, 0, 0, 0,
  1.069057e-013, 3.759135e-014, 4.089436e-011, 1.006705e-010,
  0, 0, 0, 0,
  1.015706e-013, 3.414807e-014, 4.131353e-011, 1.223027e-010,
  0, 0, 0, 0,
  4.218625e-013, 9.38207e-014, 1.462923e-010, 4.243324e-010,
  0, 0, 0, 0,
  2.672495e-013, 8.424025e-014, 1.350736e-010, 4.047384e-010,
  0, 0, 0, 0,
  1.381667e-013, 1.018631e-013, 8.926669e-011, 2.057631e-010,
  0, 0, 0, 0,
  1.103545e-013, 5.742622e-014, 6.633315e-011, 1.388415e-010,
  0, 0, 0, 0,
  2.374092e-013, 6.492612e-014, 6.687419e-011, 1.739871e-010,
  0, 0, 0, 0,
  1.104341e-013, 8.098555e-014, 5.375395e-011, 9.978517e-011,
  0, 0, 0, 0,
  1.74714e-013, 5.768629e-014, 5.504293e-011, 1.662998e-010,
  0, 0, 0, 0,
  1.644475e-013, 3.558142e-014, 6.090212e-011, 1.919095e-010,
  0, 0, 0, 0,
  9.81248e-014, 5.201194e-014, 3.396294e-011, 9.681347e-011,
  0, 0, 0, 0,
  7.758063e-014, 2.216372e-014, 2.952843e-011, 8.159182e-011,
  0, 0, 0, 0,
  1.418655e-013, 3.694661e-014, 4.984238e-011, 1.737833e-010,
  0, 0, 0, 0,
  1.182739e-013, 4.379634e-014, 3.086742e-011, 9.441502e-011,
  0, 0, 0, 0,
  5.954681e-014, 3.70309e-014, 2.959723e-011, 8.287473e-011,
  0, 0, 0, 0,
  5.829034e-014, 4.476513e-014, 4.210467e-011, 8.08935e-011,
  0, 0, 0, 0,
  3.036261e-014, 4.143692e-014, 4.408057e-011, 9.804701e-011,
  0, 0, 0, 0,
  1.094153e-013, 3.392822e-014, 3.643428e-011, 9.176846e-011,
  0, 0, 0, 0,
  5.503674e-014, 2.862366e-014, 5.196366e-011, 9.440887e-011,
  0, 0, 0, 0,
  4.684698e-014, 2.726965e-014, 2.997603e-011, 7.561424e-011,
  0, 0, 0, 0,
  1.916941e-013, 4.990986e-014, 8.309645e-011, 2.886031e-010,
  0, 0, 0, 0,
  1.089233e-013, 5.608298e-014, 4.429453e-011, 1.112334e-010,
  0, 0, 0, 0,
  1.300693e-013, 3.739233e-014, 6.725141e-011, 1.846761e-010,
  0, 0, 0, 0,
  1.73794e-013, 4.441975e-014, 5.701198e-011, 1.796391e-010,
  0, 0, 0, 0,
  6.388999e-013, 1.349722e-013, 1.801139e-010, 6.118983e-010,
  0, 0, 0, 0,
  2.345231e-013, 9.651152e-014, 1.068075e-010, 2.653964e-010,
  0, 0, 0, 0,
  1.591997e-013, 9.185172e-014, 9.540382e-011, 1.975087e-010,
  0, 0, 0, 0,
  1.507706e-013, 1.221206e-013, 1.097545e-010, 2.566777e-010,
  0, 0, 0, 0,
  1.538144e-013, 9.175175e-014, 8.688155e-011, 1.892458e-010,
  0, 0, 0, 0,
  1.097864e-013, 7.743691e-014, 6.92103e-011, 1.491144e-010,
  0, 0, 0, 0,
  7.091739e-015, 3.339166e-015, 3.157547e-012, 3.256067e-012,
  0, 0, 0, 0,
  3.294149e-014, 6.076472e-015, 4.882041e-011, 3.899402e-011,
  0, 0, 0, 0,
  1.142625e-013, 1.784391e-014, 4.721057e-012, 4.870422e-012,
  0, 0, 0, 0,
  8.092349e-015, 1.365325e-014, 8.977474e-012, 1.242688e-011,
  0, 0, 0, 0,
  5.77627e-015, 5.135203e-015, 4.723832e-012, 6.806752e-012,
  0, 0, 0, 0,
  6.290963e-015, 3.701473e-015, 1.218143e-011, 1.4051e-011,
  0, 0, 0, 0,
  9.004906e-014, 1.810883e-014, 1.066326e-011, 1.010524e-011,
  0, 0, 0, 0,
  3.94831e-015, 8.738534e-015, 8.116685e-012, 1.289421e-011,
  0, 0, 0, 0,
  6.148736e-015, 4.126315e-015, 1.457787e-011, 6.261525e-012,
  0, 0, 0, 0,
  2.957602e-014, 1.894056e-013, 1.829487e-011, 1.477625e-011,
  0, 0, 0, 0,
  8.892325e-014, 1.657996e-014, 2.464617e-012, 2.830513e-012,
  0, 0, 0, 0,
  1.088748e-014, 4.074474e-015, 3.090467e-012, 3.222225e-012,
  0, 0, 0, 0,
  3.542732e-015, 2.680905e-015, 8.498533e-012, 7.399562e-012,
  0, 0, 0, 0,
  4.826335e-015, 2.995812e-015, 3.991563e-012, 3.998955e-012,
  0, 0, 0, 0,
  3.103038e-015, 3.202749e-015, 1.721587e-012, 2.029201e-012,
  0, 0, 0, 0,
  4.050606e-015, 3.362283e-015, 4.275328e-012, 5.255847e-012,
  0, 0, 0, 0,
  5.521765e-015, 3.312049e-015, 9.528661e-012, 1.558463e-011,
  0, 0, 0, 0,
  4.155852e-015, 4.582662e-015, 2.636488e-012, 3.445081e-012,
  0, 0, 0, 0,
  4.995149e-015, 1.224269e-014, 2.719519e-012, 3.75948e-012,
  0, 0, 0, 0,
  3.990858e-015, 5.895722e-015, 4.914172e-012, 1.110442e-011,
  0, 0, 0, 0,
  2.962859e-015, 1.881475e-015, 5.500335e-012, 9.220913e-012,
  0, 0, 0, 0,
  2.884559e-015, 2.347672e-015, 3.856683e-012, 3.679512e-012,
  0, 0, 0, 0,
  1.010616e-014, 3.134504e-015, 5.095202e-012, 7.484896e-012,
  0, 0, 0, 0,
  9.017127e-014, 1.426712e-014, 7.209732e-012, 1.25441e-011,
  0, 0, 0, 0,
  5.166138e-015, 1.273123e-014, 4.257771e-012, 5.4678e-012,
  0, 0, 0, 0,
  3.652164e-015, 6.603998e-015, 1.313454e-011, 1.459086e-011,
  0, 0, 0, 0,
  5.443747e-015, 1.42385e-014, 7.357182e-012, 9.014598e-012,
  0, 0, 0, 0,
  9.594737e-014, 1.546074e-014, 1.177168e-011, 1.180514e-011,
  0, 0, 0, 0,
  4.313546e-015, 5.703668e-015, 4.969024e-012, 6.349633e-012,
  0, 0, 0, 0,
  5.13343e-015, 4.137498e-015, 4.800264e-012, 2.670465e-012,
  0, 0, 0, 0,
  3.523877e-015, 2.52465e-015, 2.674933e-012, 2.220948e-012,
  0, 0, 0, 0,
  7.868112e-015, 3.275891e-015, 8.740661e-012, 4.260821e-011,
  0, 0, 0, 0,
  4.299787e-015, 2.745928e-015, 4.487878e-012, 3.368289e-012,
  0, 0, 0, 0,
  1.852235e-014, 3.799113e-015, 1.089157e-011, 3.668207e-011,
  0, 0, 0, 0,
  8.616051e-015, 3.207253e-015, 8.552701e-012, 1.928104e-011,
  0, 0, 0, 0,
  7.690822e-014, 1.276452e-014, 6.638075e-012, 7.21721e-012,
  0, 0, 0, 0,
  9.136404e-014, 1.450296e-014, 1.173165e-011, 2.339704e-011,
  0, 0, 0, 0,
  3.688921e-015, 2.225913e-015, 2.537827e-012, 2.615865e-012,
  0, 0, 0, 0,
  3.744205e-015, 3.167416e-015, 1.527985e-012, 1.602066e-012,
  0, 0, 0, 0,
  1.552683e-014, 3.883105e-015, 2.512293e-012, 3.172591e-012,
  0, 0, 0, 0,
  7.719732e-014, 1.229547e-014, 3.212556e-012, 3.144581e-012,
  0, 0, 0, 0,
  6.218802e-015, 2.604286e-015, 7.296578e-012, 7.086357e-012,
  0, 0, 0, 0,
  2.672652e-015, 3.229974e-015, 2.494924e-012, 2.937305e-012,
  0, 0, 0, 0,
  4.1108e-015, 3.916216e-015, 2.492905e-012, 3.874205e-012,
  0, 0, 0, 0,
  9.610664e-014, 1.516244e-014, 2.065931e-012, 2.021788e-012,
  0, 0, 0, 0,
  1.321464e-014, 3.296886e-015, 2.275334e-012, 3.011622e-012,
  0, 0, 0, 0,
  6.155044e-015, 3.286652e-014, 6.225298e-012, 1.054166e-011,
  0, 0, 0, 0,
  5.79076e-015, 1.204161e-014, 2.834782e-012, 4.13132e-012,
  0, 0, 0, 0,
  1.350843e-013, 6.625909e-014, 8.519181e-012, 1.315197e-011,
  0, 0, 0, 0,
  1.793993e-014, 5.015371e-015, 1.177698e-011, 1.310601e-011,
  0, 0, 0, 0,
  4.491988e-015, 3.306506e-015, 2.239818e-012, 2.333207e-012,
  0, 0, 0, 0,
  2.79815e-015, 3.42138e-015, 2.147915e-012, 2.857288e-012,
  0, 0, 0, 0,
  5.064056e-014, 8.323637e-015, 4.554144e-012, 4.110601e-012,
  0, 0, 0, 0,
  3.742839e-014, 6.627931e-015, 5.666359e-012, 1.116606e-011,
  0, 0, 0, 0,
  3.020096e-015, 2.578346e-015, 2.275556e-012, 2.065039e-012,
  0, 0, 0, 0,
  4.036093e-015, 4.740728e-015, 2.51993e-012, 2.983695e-012,
  0, 0, 0, 0,
  2.731847e-014, 4.641794e-015, 2.824469e-012, 3.547642e-012,
  0, 0, 0, 0,
  6.835238e-014, 1.206361e-014, 3.067054e-012, 3.899706e-012,
  0, 0, 0, 0,
  2.63443e-015, 6.44804e-015, 2.366023e-012, 2.474798e-012,
  0, 0, 0, 0,
  3.984191e-015, 3.075085e-015, 1.944138e-012, 2.189714e-012,
  0, 0, 0, 0,
  2.876972e-015, 2.679468e-015, 1.960115e-012, 1.854366e-012,
  0, 0, 0, 0,
  2.26363e-015, 3.203153e-015, 1.62093e-012, 1.908999e-012,
  0, 0, 0, 0,
  3.238253e-015, 3.010812e-015, 1.959643e-012, 1.622973e-012,
  0, 0, 0, 0,
  1.848926e-015, 2.404606e-015, 1.790786e-012, 1.390343e-012,
  0, 0, 0, 0,
  2.490598e-015, 3.310425e-015, 2.481771e-012, 1.561285e-012,
  0, 0, 0, 0,
  1.377887e-013, 2.171972e-014, 3.748907e-012, 4.590315e-012,
  0, 0, 0, 0,
  5.837699e-015, 3.996839e-015, 3.412089e-012, 4.416945e-012,
  0, 0, 0, 0,
  3.964444e-015, 7.531736e-015, 8.572004e-012, 1.236402e-011,
  0, 0, 0, 0,
  4.884795e-015, 8.160531e-015, 1.145919e-011, 1.497409e-011,
  0, 0, 0, 0,
  6.761499e-014, 1.086004e-014, 6.396136e-012, 1.151573e-011,
  0, 0, 0, 0,
  2.023375e-014, 3.859621e-015, 3.862132e-012, 3.844641e-012,
  0, 0, 0, 0,
  4.427194e-015, 4.352518e-015, 1.235501e-011, 1.396292e-011,
  0, 0, 0, 0,
  4.171055e-015, 2.711501e-015, 2.850827e-012, 4.255778e-012,
  0, 0, 0, 0,
  3.816151e-014, 7.076099e-015, 2.428013e-012, 3.005154e-012,
  0, 0, 0, 0,
  5.60485e-014, 8.978147e-015, 2.825288e-012, 2.145257e-012,
  0, 0, 0, 0,
  4.621567e-015, 3.418192e-015, 3.769155e-012, 3.224196e-012,
  0, 0, 0, 0,
  7.521249e-015, 3.452332e-015, 1.872853e-012, 1.878703e-012,
  0, 0, 0, 0,
  9.673631e-015, 4.754706e-015, 4.428566e-012, 4.940209e-012,
  0, 0, 0, 0,
  6.420296e-015, 4.006454e-015, 8.720079e-012, 1.117862e-011,
  0, 0, 0, 0,
  4.996614e-015, 5.607823e-015, 3.805975e-012, 6.241371e-012,
  0, 0, 0, 0,
  4.955456e-015, 6.692044e-015, 4.020151e-012, 5.834967e-012,
  0, 0, 0, 0,
  3.433968e-015, 5.487193e-015, 7.235687e-012, 1.044157e-011,
  0, 0, 0, 0,
  1.521206e-013, 2.376647e-014, 6.451877e-012, 8.187247e-012,
  0, 0, 0, 0,
  5.835454e-015, 1.249517e-014, 9.875837e-012, 2.378997e-011,
  0, 0, 0, 0,
  7.107109e-015, 5.72954e-015, 8.417193e-012, 1.084821e-011,
  0, 0, 0, 0,
  5.170233e-015, 5.839316e-015, 5.698005e-012, 8.272394e-012,
  0, 0, 0, 0,
  8.063992e-014, 1.299645e-014, 5.170244e-012, 5.123366e-012,
  0, 0, 0, 0,
  1.140528e-014, 5.738483e-015, 4.388157e-012, 7.712973e-012,
  0, 0, 0, 0,
  5.070254e-015, 3.685575e-015, 7.088283e-012, 9.269484e-012,
  0, 0, 0, 0,
  5.77905e-015, 1.703814e-014, 1.406934e-011, 2.284047e-011,
  0, 0, 0, 0,
  6.071716e-014, 1.394389e-014, 1.177123e-011, 2.063933e-011,
  0, 0, 0, 0,
  3.632321e-014, 8.090046e-015, 4.386018e-012, 6.951285e-012,
  0, 0, 0, 0,
  5.558591e-015, 1.352987e-014, 9.163838e-012, 8.900666e-012,
  0, 0, 0, 0,
  1.765358e-014, 5.22987e-015, 1.387401e-011, 1.445785e-011,
  0, 0, 0, 0,
  2.621442e-014, 1.979343e-014, 1.241364e-011, 2.729739e-011,
  0, 0, 0, 0,
  3.277141e-015, 2.736252e-015, 4.742067e-012, 5.980107e-012,
  0, 0, 0, 0,
  3.342744e-015, 2.394366e-015, 4.205749e-012, 4.037157e-012,
  0, 0, 0, 0,
  8.086281e-015, 4.145083e-015, 2.968934e-012, 4.862064e-012,
  0, 0, 0, 0,
  4.243972e-015, 5.120027e-015, 6.240279e-012, 7.650495e-012,
  0, 0, 0, 0,
  6.073325e-015, 4.147974e-015, 1.863437e-012, 1.635462e-012,
  0, 0, 0, 0,
  4.026855e-015, 3.013802e-015, 1.401606e-012, 1.488112e-012,
  0, 0, 0, 0,
  7.772634e-015, 6.380356e-015, 1.986425e-012, 2.049109e-012,
  0, 0, 0, 0,
  8.259122e-014, 1.332829e-014, 1.080516e-011, 1.904037e-011,
  0, 0, 0, 0,
  4.113971e-014, 7.888808e-015, 7.627499e-011, 8.275953e-011,
  0, 0, 0, 0,
  1.539245e-014, 9.618187e-015, 4.772582e-011, 5.603045e-011,
  0, 0, 0, 0,
  8.616216e-014, 2.495326e-014, 2.187275e-011, 3.363718e-011,
  0, 0, 0, 0,
  8.876485e-015, 4.980573e-015, 5.65674e-012, 7.079729e-012,
  0, 0, 0, 0,
  1.015674e-014, 7.305612e-015, 5.130823e-012, 9.581682e-012,
  0, 0, 0, 0,
  1.453256e-014, 1.552822e-014, 1.77739e-011, 2.977192e-011,
  0, 0, 0, 0,
  1.351509e-014, 5.954829e-015, 5.250607e-012, 1.010521e-011,
  0, 0, 0, 0,
  8.909372e-015, 4.98891e-015, 5.871002e-012, 7.975243e-012,
  0, 0, 0, 0,
  1.240854e-014, 4.468844e-015, 3.135725e-012, 7.182858e-012,
  0, 0, 0, 0,
  1.075491e-014, 6.007403e-015, 3.550573e-012, 7.580633e-012,
  0, 0, 0, 0,
  2.72063e-014, 6.933446e-015, 5.684985e-012, 1.16588e-011,
  0, 0, 0, 0,
  4.478494e-014, 9.486412e-015, 1.660636e-011, 3.304217e-011,
  0, 0, 0, 0,
  4.719103e-014, 9.88259e-015, 1.797383e-011, 2.60178e-011,
  0, 0, 0, 0,
  3.94017e-014, 9.535497e-015, 4.155688e-012, 8.572831e-012,
  0, 0, 0, 0,
  6.095677e-014, 1.826756e-014, 6.08056e-012, 1.460131e-011,
  0, 0, 0, 0,
  1.726919e-013, 3.882727e-014, 5.940424e-012, 3.0719e-011,
  0, 0, 0, 0,
  4.541684e-013, 7.686456e-014, 1.186748e-011, 4.033333e-011,
  0, 0, 0, 0,
  3.591882e-013, 6.953684e-014, 7.870573e-012, 3.765342e-011,
  0, 0, 0, 0,
  8.552929e-013, 1.542017e-013, 2.367125e-011, 1.002535e-010,
  0, 0, 0, 0,
  7.310108e-013, 1.444634e-013, 1.879369e-011, 6.131484e-011,
  0, 0, 0, 0,
  1.891734e-012, 3.759587e-013, 6.106161e-011, 2.687643e-010,
  0, 0, 0, 0,
  2.695332e-012, 5.289674e-013, 1.432882e-010, 4.741454e-010,
  0, 0, 0, 0,
  2.799352e-012, 8.211796e-013, 1.105902e-010, 4.173627e-010,
  0, 0, 0, 0,
  4.469326e-012, 1.044354e-012, 2.032637e-010, 8.02687e-010,
  0, 0, 0, 0,
  1.129483e-011, 2.890218e-012, 7.713706e-010, 2.326421e-009,
  0, 0, 0, 0,
  1.70495e-011, 4.844641e-012, 1.545121e-009, 7.682195e-009,
  0, 0, 0, 0,
  2.363355e-011, 6.48167e-012, 1.486892e-009, 5.514919e-009,
  0, 0, 0, 0,
  1.801467e-011, 5.298257e-012, 1.348143e-009, 4.857211e-009,
  0, 0, 0, 0,
  1.576294e-011, 5.436223e-012, 1.203013e-009, 3.956691e-009,
  0, 0, 0, 0,
  1.663664e-011, 6.777877e-012, 1.447625e-009, 5.969226e-009,
  0, 0, 0, 0,
  6.014823e-012, 2.389909e-012, 4.263799e-010, 1.687859e-009,
  0, 0, 0, 0,
  4.1162e-012, 7.735028e-013, 1.575415e-010, 6.763066e-010,
  0, 0, 0, 0,
  2.2183e-012, 6.024098e-013, 8.042945e-011, 3.407002e-010,
  0, 0, 0, 0,
  2.113684e-012, 5.411394e-013, 7.117586e-011, 3.247816e-010,
  0, 0, 0, 0,
  9.345819e-013, 3.8495e-013, 8.769951e-011, 1.445492e-010,
  0, 0, 0, 0,
  5.933906e-013, 5.103276e-013, 1.431685e-010, 2.873812e-010,
  0, 0, 0, 0,
  3.638419e-013, 4.185538e-013, 5.192683e-011, 1.161217e-010,
  0, 0, 0, 0,
  5.177425e-013, 4.134206e-013, 2.743833e-011, 5.59259e-011,
  0, 0, 0, 0,
  3.062539e-013, 1.017526e-013, 2.485193e-011, 5.216633e-011,
  0, 0, 0, 0,
  2.087113e-013, 7.685816e-014, 4.458737e-011, 9.659622e-011,
  0, 0, 0, 0,
  7.29769e-014, 5.367914e-014, 3.369117e-011, 7.21365e-011,
  0, 0, 0, 0,
  1.18667e-013, 2.920004e-014, 1.565717e-011, 3.550106e-011,
  0, 0, 0, 0,
  5.816007e-014, 1.329876e-013, 1.05599e-010, 2.364053e-010,
  0, 0, 0, 0,
  3.040609e-014, 1.161542e-014, 1.16705e-011, 2.146115e-011,
  0, 0, 0, 0,
  2.087757e-014, 1.499416e-014, 1.168958e-011, 2.277457e-011,
  0, 0, 0, 0,
  1.336155e-014, 2.166016e-014, 1.678601e-011, 3.618652e-011,
  0, 0, 0, 0,
  2.290818e-014, 1.444279e-014, 1.285101e-011, 2.253689e-011,
  0, 0, 0, 0,
  2.736299e-014, 1.257997e-013, 7.309942e-011, 1.62444e-010,
  0, 0, 0, 0,
  3.042655e-014, 1.758253e-013, 1.243e-010, 2.713731e-010,
  0, 0, 0, 0,
  4.148329e-014, 2.387005e-013, 2.666314e-010, 6.310219e-010,
  0, 0, 0, 0,
  9.751655e-014, 3.287061e-013, 2.02856e-010, 4.315384e-010,
  0, 0, 0, 0,
  3.476866e-014, 2.140003e-013, 1.399019e-010, 3.054688e-010,
  0, 0, 0, 0,
  3.356417e-014, 2.122841e-013, 1.652039e-010, 3.581742e-010,
  0, 0, 0, 0,
  1.19516e-014, 3.249494e-014, 2.455845e-011, 5.816566e-011,
  0, 0, 0, 0,
  1.41159e-014, 7.774041e-014, 6.031531e-011, 1.326354e-010,
  0, 0, 0, 0,
  1.154127e-014, 6.337704e-014, 3.966144e-011, 9.398432e-011,
  0, 0, 0, 0,
  7.19289e-015, 4.842963e-015, 1.281804e-011, 1.319967e-011,
  0, 0, 0, 0,
  4.345543e-015, 5.868223e-015, 5.655626e-012, 7.458502e-012,
  0, 0, 0, 0,
  5.16572e-015, 2.590587e-014, 1.666332e-011, 3.258136e-011,
  0, 0, 0, 0,
  4.338009e-015, 9.282725e-015, 6.499081e-012, 1.273141e-011,
  0, 0, 0, 0,
  5.893907e-015, 7.514448e-015, 5.458918e-012, 8.962528e-012,
  0, 0, 0, 0,
  4.0528e-015, 1.154209e-014, 8.761659e-012, 1.723172e-011,
  0, 0, 0, 0,
  3.148908e-014, 2.827361e-014, 2.252268e-011, 5.575826e-011,
  0, 0, 0, 0,
  6.481348e-015, 1.808599e-014, 1.549232e-011, 3.543226e-011,
  0, 0, 0, 0,
  2.570677e-014, 1.629691e-013, 1.202152e-010, 2.730549e-010,
  0, 0, 0, 0,
  4.509898e-014, 2.880695e-013, 2.099957e-010, 4.786894e-010,
  0, 0, 0, 0,
  1.422491e-013, 9.251552e-013, 4.229147e-010, 9.330076e-010,
  0, 0, 0, 0,
  1.469549e-013, 1.833962e-013, 1.176299e-010, 2.644176e-010,
  0, 0, 0, 0,
  3.994316e-014, 2.58162e-013, 1.518204e-010, 3.299465e-010,
  0, 0, 0, 0,
  2.51454e-014, 1.589008e-013, 1.187968e-010, 2.695104e-010,
  0, 0, 0, 0,
  1.863636e-014, 1.138708e-013, 8.093538e-011, 1.889697e-010,
  0, 0, 0, 0,
  7.505894e-014, 1.072617e-013, 7.906105e-011, 1.968953e-010,
  0, 0, 0, 0,
  3.185184e-014, 1.902725e-013, 1.45981e-010, 3.35398e-010,
  0, 0, 0, 0,
  7.786798e-015, 4.325648e-014, 3.015197e-011, 7.357852e-011,
  0, 0, 0, 0,
  9.4405e-015, 4.557022e-014, 3.025602e-011, 7.39209e-011,
  0, 0, 0, 0,
  6.390912e-014, 2.089684e-013, 1.458007e-010, 3.342512e-010,
  0, 0, 0, 0,
  3.570702e-014, 5.65303e-014, 4.437036e-011, 9.584145e-011,
  0, 0, 0, 0,
  3.96668e-014, 2.517581e-013, 1.948583e-010, 4.405932e-010,
  0, 0, 0, 0,
  1.145991e-014, 5.38294e-014, 4.450981e-011, 9.313812e-011,
  0, 0, 0, 0,
  1.890038e-014, 7.634811e-014, 8.701612e-011, 1.740621e-010,
  0, 0, 0, 0,
  3.820224e-014, 1.553213e-013, 1.110507e-010, 2.572185e-010,
  0, 0, 0, 0,
  4.292786e-014, 2.774395e-013, 1.84876e-010, 4.07332e-010,
  0, 0, 0, 0,
  2.992127e-014, 1.891146e-013, 1.571531e-010, 3.544766e-010,
  0, 0, 0, 0,
  8.318675e-014, 5.391252e-013, 2.933213e-010, 6.849574e-010,
  0, 0, 0, 0,
  1.404095e-013, 2.138403e-013, 1.561833e-010, 3.592573e-010,
  0, 0, 0, 0,
  7.841021e-014, 5.092733e-013, 3.594848e-010, 8.088948e-010,
  0, 0, 0, 0,
  4.858656e-014, 3.117165e-013, 2.3217e-010, 5.357121e-010,
  0, 0, 0, 0,
  5.967384e-014, 3.852781e-013, 2.702799e-010, 6.214927e-010,
  0, 0, 0, 0,
  8.137925e-014, 2.903843e-014, 1.185829e-011, 2.503495e-011,
  0, 0, 0, 0,
  1.039199e-014, 5.832809e-014, 4.206974e-011, 9.837312e-011,
  0, 0, 0, 0,
  1.899891e-014, 1.168829e-013, 8.564959e-011, 2.014245e-010,
  0, 0, 0, 0,
  1.222719e-014, 6.715047e-014, 4.585974e-011, 1.104593e-010,
  0, 0, 0, 0,
  6.712578e-014, 3.009123e-014, 2.474076e-011, 5.341645e-011,
  0, 0, 0, 0,
  2.30388e-014, 7.779164e-015, 7.175916e-012, 1.208546e-011,
  0, 0, 0, 0,
  3.483118e-015, 9.157308e-015, 1.069392e-011, 1.606327e-011,
  0, 0, 0, 0,
  4.529277e-015, 7.51737e-015, 7.262803e-012, 1.042095e-011,
  0, 0, 0, 0,
  1.613501e-014, 9.665527e-014, 7.006053e-011, 1.634097e-010,
  0, 0, 0, 0,
  2.135076e-014, 1.353092e-013, 1.00949e-010, 2.354312e-010,
  0, 0, 0, 0,
  1.121536e-014, 6.992554e-014, 4.750929e-011, 1.104862e-010,
  0, 0, 0, 0,
  1.625543e-014, 1.023718e-013, 7.31105e-011, 1.65651e-010,
  0, 0, 0, 0,
  2.683192e-014, 4.784775e-014, 4.348203e-011, 8.718547e-011,
  0, 0, 0, 0,
  1.442063e-013, 1.05147e-013, 6.747328e-011, 1.525642e-010,
  0, 0, 0, 0,
  2.256553e-014, 1.447219e-013, 1.237287e-010, 2.790281e-010,
  0, 0, 0, 0,
  7.569959e-014, 3.732744e-013, 2.689141e-010, 5.931431e-010,
  0, 0, 0, 0,
  1.591202e-013, 2.479407e-013, 2.272668e-010, 5.775002e-010,
  0, 0, 0, 0,
  1.054031e-013, 4.076267e-013, 3.303095e-010, 7.42565e-010,
  0, 0, 0, 0,
  1.105004e-013, 6.532678e-013, 5.25215e-010, 1.18528e-009,
  0, 0, 0, 0,
  3.214468e-013, 3.928591e-013, 2.142237e-010, 5.61533e-010,
  0, 0, 0, 0,
  1.232001e-013, 3.749567e-013, 2.717446e-010, 6.173397e-010,
  0, 0, 0, 0,
  1.73885e-013, 2.824813e-013, 2.36561e-010, 5.601682e-010,
  0, 0, 0, 0,
  1.067814e-013, 1.241678e-013, 1.556897e-010, 3.841638e-010,
  0, 0, 0, 0,
  3.808907e-013, 9.931062e-014, 2.220653e-010, 7.4422e-010,
  0, 0, 0, 0,
  1.713299e-013, 9.786429e-014, 1.111319e-010, 3.438844e-010,
  0, 0, 0, 0,
  4.77968e-013, 1.758334e-013, 2.202066e-010, 7.763961e-010,
  0, 0, 0, 0,
  1.799784e-013, 7.662374e-014, 1.342922e-010, 4.301997e-010,
  0, 0, 0, 0,
  7.12005e-013, 1.77259e-013, 3.384057e-010, 1.236043e-009,
  0, 0, 0, 0,
  3.433322e-013, 1.978768e-013, 3.213255e-010, 9.180706e-010,
  0, 0, 0, 0,
  9.609177e-014, 1.01773e-013, 1.160394e-010, 3.16459e-010,
  0, 0, 0, 0,
  1.486627e-013, 8.813739e-014, 9.495381e-011, 2.823917e-010,
  0, 0, 0, 0,
  2.239761e-013, 1.620763e-013, 1.036337e-010, 3.184327e-010,
  0, 0, 0, 0,
  2.594901e-014, 2.413239e-014, 3.457046e-011, 6.65289e-011,
  0, 0, 0, 0,
  2.489202e-014, 3.821935e-014, 3.483327e-011, 8.700763e-011,
  0, 0, 0, 0,
  8.589651e-014, 9.772046e-014, 8.512446e-011, 2.229639e-010,
  0, 0, 0, 0,
  1.97e-014, 7.612667e-014, 6.141478e-011, 1.439764e-010,
  0, 0, 0, 0,
  9.413037e-015, 4.692945e-015, 5.929101e-012, 1.653965e-011,
  0, 0, 0, 0,
  1.170449e-014, 4.21011e-015, 8.628992e-012, 1.777601e-011,
  0, 0, 0, 0,
  4.277849e-015, 7.916738e-015, 5.568771e-012, 1.476099e-011,
  0, 0, 0, 0,
  4.89555e-015, 6.083219e-015, 5.051332e-012, 8.47352e-012,
  0, 0, 0, 0,
  4.959037e-015, 3.399334e-015, 8.772004e-012, 1.128668e-011,
  0, 0, 0, 0,
  1.381797e-014, 8.905626e-015, 7.282206e-012, 1.243056e-011,
  0, 0, 0, 0,
  5.956233e-014, 1.851718e-014, 1.70641e-011, 3.681803e-011,
  0, 0, 0, 0,
  2.854417e-014, 5.220291e-014, 4.362239e-011, 9.551964e-011,
  0, 0, 0, 0,
  1.60086e-014, 9.377637e-014, 6.742896e-011, 1.634072e-010,
  0, 0, 0, 0,
  7.781693e-015, 3.562461e-014, 2.727146e-011, 6.32813e-011,
  0, 0, 0, 0,
  3.067876e-014, 1.090449e-014, 1.239604e-011, 2.390643e-011,
  0, 0, 0, 0,
  7.666118e-014, 2.768654e-014, 2.765575e-011, 9.060443e-011,
  0, 0, 0, 0,
  2.804567e-013, 4.693903e-014, 1.425598e-010, 4.982148e-010,
  0, 0, 0, 0,
  8.812301e-014, 2.255972e-014, 7.894384e-011, 2.335442e-010,
  0, 0, 0, 0,
  1.192293e-013, 2.63134e-014, 6.809144e-011, 2.247659e-010,
  0, 0, 0, 0,
  4.347388e-013, 1.269442e-013, 2.307405e-010, 7.506299e-010,
  0, 0, 0, 0,
  3.137081e-013, 4.891316e-014, 1.619356e-010, 5.488329e-010,
  0, 0, 0, 0,
  2.365288e-013, 3.669278e-014, 1.214812e-010, 4.139632e-010,
  0, 0, 0, 0,
  4.998016e-013, 7.883344e-014, 2.727777e-010, 9.239903e-010,
  0, 0, 0, 0,
  4.57805e-013, 7.113058e-014, 2.094621e-010, 7.583866e-010,
  0, 0, 0, 0,
  1.107339e-013, 4.431662e-014, 9.384486e-011, 2.682652e-010,
  0, 0, 0, 0,
  1.589257e-013, 1.667862e-013, 2.031805e-010, 5.732202e-010,
  0, 0, 0, 0,
  4.513597e-013, 1.00499e-013, 2.793672e-010, 9.592996e-010,
  0, 0, 0, 0,
  3.835892e-013, 2.441811e-013, 3.397578e-010, 9.117818e-010,
  0, 0, 0, 0,
  6.58346e-013, 4.010045e-013, 4.867636e-010, 1.426494e-009,
  0, 0, 0, 0,
  5.396797e-013, 3.127591e-013, 3.082298e-010, 9.829343e-010,
  0, 0, 0, 0,
  4.888504e-013, 3.539784e-013, 2.720871e-010, 7.360322e-010,
  0, 0, 0, 0,
  8.087205e-013, 2.776356e-013, 3.804276e-010, 1.196236e-009,
  0, 0, 0, 0,
  5.303242e-013, 1.919938e-013, 4.06207e-010, 1.265567e-009,
  0, 0, 0, 0,
  1.647125e-013, 5.981944e-014, 1.017942e-010, 3.251152e-010,
  0, 0, 0, 0,
  6.622606e-014, 3.394531e-014, 5.541002e-011, 1.428422e-010,
  0, 0, 0, 0,
  2.641019e-013, 4.746624e-014, 1.425659e-010, 4.935831e-010,
  0, 0, 0, 0,
  8.651136e-014, 1.573251e-014, 2.169466e-011, 6.105265e-011,
  0, 0, 0, 0,
  2.640782e-014, 1.269753e-014, 1.900769e-011, 4.912361e-011,
  0, 0, 0, 0,
  1.595467e-014, 1.262893e-014, 1.543846e-011, 2.673175e-011,
  0, 0, 0, 0,
  1.317683e-014, 9.404492e-015, 2.079926e-011, 2.672594e-011,
  0, 0, 0, 0,
  9.931086e-014, 1.630222e-014, 1.519529e-011, 4.222341e-011,
  0, 0, 0, 0,
  1.339971e-014, 1.539031e-014, 1.339621e-011, 2.310666e-011,
  0, 0, 0, 0,
  2.335428e-013, 1.593898e-013, 1.401397e-010, 4.13052e-010,
  0, 0, 0, 0,
  2.244055e-013, 3.603587e-013, 1.759976e-010, 4.250074e-010,
  0, 0, 0, 0,
  5.563605e-014, 1.320358e-013, 1.237399e-010, 2.927479e-010,
  0, 0, 0, 0,
  8.069154e-014, 1.357889e-013, 1.352738e-010, 3.264212e-010,
  0, 0, 0, 0,
  8.332029e-014, 1.94947e-013, 1.496146e-010, 3.506966e-010,
  0, 0, 0, 0,
  3.184422e-013, 1.675291e-013, 1.858632e-010, 6.008395e-010,
  0, 0, 0, 0,
  2.822809e-013, 1.900727e-013, 2.182555e-010, 6.224305e-010,
  0, 0, 0, 0,
  4.00461e-013, 1.077098e-013, 2.23149e-010, 7.456379e-010,
  0, 0, 0, 0,
  3.837962e-013, 9.737764e-014, 2.366442e-010, 7.897824e-010,
  0, 0, 0, 0,
  4.754046e-014, 1.021918e-013, 9.137858e-011, 2.100423e-010,
  0, 0, 0, 0,
  3.384498e-013, 9.220638e-014, 2.228046e-010, 7.007951e-010,
  0, 0, 0, 0,
  7.232552e-013, 1.219576e-013, 3.562179e-010, 1.228188e-009,
  0, 0, 0, 0,
  3.064497e-013, 1.052272e-013, 2.102884e-010, 6.378829e-010,
  0, 0, 0, 0,
  2.593324e-013, 6.458723e-014, 1.449091e-010, 4.950757e-010,
  0, 0, 0, 0,
  2.192831e-013, 6.509771e-014, 1.137236e-010, 3.896648e-010,
  0, 0, 0, 0,
  8.569896e-014, 6.201576e-014, 5.860626e-011, 1.387413e-010,
  0, 0, 0, 0,
  3.129019e-014, 2.611415e-014, 2.959425e-011, 8.529898e-011,
  0, 0, 0, 0,
  7.635878e-014, 8.656946e-014, 6.913176e-011, 1.942255e-010,
  0, 0, 0, 0,
  2.426914e-013, 4.619774e-014, 1.267861e-010, 4.209205e-010,
  0, 0, 0, 0,
  1.18657e-013, 1.56459e-013, 1.0721e-010, 3.113301e-010,
  0, 0, 0, 0,
  7.37991e-014, 3.493441e-014, 5.749468e-011, 1.575038e-010,
  0, 0, 0, 0,
  3.524014e-013, 5.856162e-014, 2.067813e-010, 6.970338e-010,
  0, 0, 0, 0,
  8.708348e-014, 5.924281e-014, 6.103896e-011, 1.935294e-010,
  0, 0, 0, 0,
  5.829768e-014, 1.350997e-013, 1.03931e-010, 2.723372e-010,
  0, 0, 0, 0,
  4.180825e-013, 9.110559e-014, 2.314244e-010, 8.035943e-010,
  0, 0, 0, 0,
  9.817278e-013, 2.695289e-013, 4.504679e-010, 1.604208e-009,
  0, 0, 0, 0,
  1.318346e-012, 3.390528e-013, 7.529554e-010, 2.511241e-009,
  0, 0, 0, 0,
  7.566373e-013, 2.654855e-013, 3.978799e-010, 1.383301e-009,
  0, 0, 0, 0,
  5.148607e-013, 2.4475e-013, 3.175968e-010, 1.029768e-009,
  0, 0, 0, 0,
  9.041355e-013, 1.589945e-013, 3.671655e-010, 1.398104e-009,
  0, 0, 0, 0,
  3.352362e-013, 2.688773e-013, 2.869999e-010, 7.601502e-010,
  0, 0, 0, 0,
  8.934225e-013, 1.962195e-013, 4.823862e-010, 1.705916e-009,
  0, 0, 0, 0,
  7.684951e-013, 1.26735e-013, 3.766455e-010, 1.391087e-009,
  0, 0, 0, 0,
  4.930264e-013, 1.138427e-013, 3.143499e-010, 1.058149e-009,
  0, 0, 0, 0,
  3.600174e-013, 6.087944e-014, 1.482256e-010, 5.789147e-010,
  0, 0, 0, 0,
  2.2236e-013, 1.002164e-013, 1.123226e-010, 3.844335e-010,
  0, 0, 0, 0,
  1.366558e-013, 3.436158e-014, 5.626243e-011, 1.905994e-010,
  0, 0, 0, 0,
  9.451151e-014, 4.092101e-014, 7.5689e-011, 2.139962e-010,
  0, 0, 0, 0,
  1.07658e-013, 1.096052e-013, 9.429642e-011, 2.487432e-010,
  0, 0, 0, 0,
  1.733031e-013, 1.088673e-013, 1.664782e-010, 4.987394e-010,
  0, 0, 0, 0,
  2.399384e-013, 1.454571e-013, 1.561711e-010, 4.963289e-010,
  0, 0, 0, 0,
  5.974978e-014, 2.355629e-014, 4.61555e-011, 1.15719e-010,
  0, 0, 0, 0,
  1.12497e-013, 3.748638e-014, 4.191259e-011, 1.535036e-010,
  0, 0, 0, 0,
  5.536482e-013, 9.064938e-014, 2.810978e-010, 1.037053e-009,
  0, 0, 0, 0,
  3.760135e-013, 1.250417e-013, 2.733231e-010, 8.505527e-010,
  0, 0, 0, 0,
  6.498089e-013, 1.176334e-013, 3.391378e-010, 1.188947e-009,
  0, 0, 0, 0,
  6.417296e-013, 1.337814e-013, 3.115835e-010, 1.131886e-009,
  0, 0, 0, 0,
  1.425196e-012, 2.761616e-013, 5.953508e-010, 2.224292e-009,
  0, 0, 0, 0,
  9.03558e-013, 4.466201e-013, 6.131426e-010, 1.94823e-009,
  0, 0, 0, 0,
  9.444758e-013, 2.679463e-013, 4.43104e-010, 1.637178e-009,
  0, 0, 0, 0,
  7.541977e-013, 2.667294e-013, 4.747695e-010, 1.467997e-009,
  0, 0, 0, 0,
  1.021172e-012, 2.959223e-013, 4.308539e-010, 1.58584e-009,
  0, 0, 0, 0,
  4.2895e-013, 2.758841e-013, 3.424274e-010, 1.025822e-009,
  0, 0, 0, 0 ;

 emf_mask =
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1,
  1, 1, 1, 1 ;
}
